
module PC ( clk, rst, PCin, PCout );
  input [31:0] PCin;
  output [31:0] PCout;
  input clk, rst;
  wire   n1, n2;

  DFFRX1 \PCout_reg[31]  ( .D(PCin[31]), .CK(clk), .RN(n1), .Q(PCout[31]) );
  DFFRX1 \PCout_reg[30]  ( .D(PCin[30]), .CK(clk), .RN(n1), .Q(PCout[30]) );
  DFFRX1 \PCout_reg[29]  ( .D(PCin[29]), .CK(clk), .RN(n1), .Q(PCout[29]) );
  DFFRX1 \PCout_reg[28]  ( .D(PCin[28]), .CK(clk), .RN(n1), .Q(PCout[28]) );
  DFFRX1 \PCout_reg[27]  ( .D(PCin[27]), .CK(clk), .RN(n1), .Q(PCout[27]) );
  DFFRX1 \PCout_reg[26]  ( .D(PCin[26]), .CK(clk), .RN(n1), .Q(PCout[26]) );
  DFFRX1 \PCout_reg[25]  ( .D(PCin[25]), .CK(clk), .RN(n1), .Q(PCout[25]) );
  DFFRX1 \PCout_reg[0]  ( .D(PCin[0]), .CK(clk), .RN(n2), .Q(PCout[0]) );
  DFFRX1 \PCout_reg[12]  ( .D(PCin[12]), .CK(clk), .RN(n2), .Q(PCout[12]) );
  DFFRX1 \PCout_reg[11]  ( .D(PCin[11]), .CK(clk), .RN(n2), .Q(PCout[11]) );
  DFFRX1 \PCout_reg[10]  ( .D(PCin[10]), .CK(clk), .RN(n2), .Q(PCout[10]) );
  DFFRX1 \PCout_reg[14]  ( .D(PCin[14]), .CK(clk), .RN(n2), .Q(PCout[14]) );
  DFFRX1 \PCout_reg[13]  ( .D(PCin[13]), .CK(clk), .RN(n2), .Q(PCout[13]) );
  DFFRX1 \PCout_reg[8]  ( .D(PCin[8]), .CK(clk), .RN(n2), .Q(PCout[8]) );
  DFFRX1 \PCout_reg[7]  ( .D(PCin[7]), .CK(clk), .RN(n2), .Q(PCout[7]) );
  DFFRX1 \PCout_reg[6]  ( .D(PCin[6]), .CK(clk), .RN(n2), .Q(PCout[6]) );
  DFFRX1 \PCout_reg[5]  ( .D(PCin[5]), .CK(clk), .RN(n2), .Q(PCout[5]) );
  DFFRX1 \PCout_reg[4]  ( .D(PCin[4]), .CK(clk), .RN(n2), .Q(PCout[4]) );
  DFFRX1 \PCout_reg[3]  ( .D(PCin[3]), .CK(clk), .RN(n2), .Q(PCout[3]) );
  DFFRX1 \PCout_reg[9]  ( .D(PCin[9]), .CK(clk), .RN(n2), .Q(PCout[9]) );
  DFFRX1 \PCout_reg[17]  ( .D(PCin[17]), .CK(clk), .RN(n2), .Q(PCout[17]) );
  DFFRX1 \PCout_reg[16]  ( .D(PCin[16]), .CK(clk), .RN(n2), .Q(PCout[16]) );
  DFFRX1 \PCout_reg[15]  ( .D(PCin[15]), .CK(clk), .RN(n2), .Q(PCout[15]) );
  DFFRX1 \PCout_reg[2]  ( .D(PCin[2]), .CK(clk), .RN(n2), .Q(PCout[2]) );
  DFFRX1 \PCout_reg[1]  ( .D(PCin[1]), .CK(clk), .RN(n2), .Q(PCout[1]) );
  DFFRX1 \PCout_reg[18]  ( .D(PCin[18]), .CK(clk), .RN(n2), .Q(PCout[18]) );
  DFFRX1 \PCout_reg[19]  ( .D(PCin[19]), .CK(clk), .RN(n2), .Q(PCout[19]) );
  DFFRX1 \PCout_reg[20]  ( .D(PCin[20]), .CK(clk), .RN(n2), .Q(PCout[20]) );
  DFFRX1 \PCout_reg[21]  ( .D(PCin[21]), .CK(clk), .RN(n2), .Q(PCout[21]) );
  DFFRX1 \PCout_reg[22]  ( .D(PCin[22]), .CK(clk), .RN(n2), .Q(PCout[22]) );
  DFFRX1 \PCout_reg[23]  ( .D(PCin[23]), .CK(clk), .RN(n2), .Q(PCout[23]) );
  DFFRX1 \PCout_reg[24]  ( .D(PCin[24]), .CK(clk), .RN(n2), .Q(PCout[24]) );
  INVX3 U3 ( .A(rst), .Y(n2) );
  CLKBUFX3 U4 ( .A(n2), .Y(n1) );
endmodule


module mainControl ( opcode_i, funct_i, RegDst_o, Jump_o, Branch_o, MemRead_o, 
        MemToReg_o, ALUOp_o, MemWrite_o, ALUSrc_o, RegWrite_o, JumpRegister_o, 
        JumpAndLink_o, Port42 );
  input [5:0] opcode_i;
  input [5:0] funct_i;
  output [1:0] ALUOp_o;
  output RegDst_o, Jump_o, Branch_o, MemRead_o, MemToReg_o, MemWrite_o,
         ALUSrc_o, RegWrite_o, JumpRegister_o, JumpAndLink_o;
  inout Port42;
  wire   n6, n7, n8, n9, n10, n11, n12, n4, n5, n13;

  CLKINVX1 U1 ( .A(n6), .Y(MemRead_o) );
  NAND3BX1 U2 ( .AN(JumpAndLink_o), .B(n6), .C(n4), .Y(RegWrite_o) );
  CLKINVX1 U3 ( .A(RegDst_o), .Y(n4) );
  NOR3X1 U4 ( .A(n13), .B(n8), .C(n5), .Y(n10) );
  CLKINVX1 U5 ( .A(n7), .Y(MemWrite_o) );
  NAND2X1 U6 ( .A(n7), .B(n6), .Y(ALUSrc_o) );
  NOR4X1 U7 ( .A(n8), .B(opcode_i[0]), .C(opcode_i[1]), .D(opcode_i[5]), .Y(
        RegDst_o) );
  NOR3X1 U8 ( .A(opcode_i[3]), .B(opcode_i[5]), .C(opcode_i[4]), .Y(n12) );
  NOR2BX1 U9 ( .AN(n10), .B(opcode_i[5]), .Y(JumpAndLink_o) );
  NAND4X1 U10 ( .A(opcode_i[5]), .B(opcode_i[1]), .C(opcode_i[3]), .D(n11), 
        .Y(n7) );
  NOR3X1 U11 ( .A(n13), .B(opcode_i[4]), .C(opcode_i[2]), .Y(n11) );
  OR3X2 U12 ( .A(opcode_i[3]), .B(opcode_i[4]), .C(opcode_i[2]), .Y(n8) );
  NAND2X1 U13 ( .A(opcode_i[5]), .B(n10), .Y(n6) );
  CLKINVX1 U14 ( .A(opcode_i[0]), .Y(n13) );
  CLKINVX1 U15 ( .A(opcode_i[1]), .Y(n5) );
  NOR4BX1 U16 ( .AN(funct_i[3]), .B(n9), .C(funct_i[0]), .D(n4), .Y(
        JumpRegister_o) );
  OR4X1 U17 ( .A(funct_i[2]), .B(funct_i[1]), .C(funct_i[5]), .D(funct_i[4]), 
        .Y(n9) );
  NOR3X1 U18 ( .A(n5), .B(opcode_i[5]), .C(n8), .Y(Jump_o) );
  CLKBUFX3 U19 ( .A(RegDst_o), .Y(ALUOp_o[1]) );
  CLKBUFX3 U20 ( .A(Branch_o), .Y(ALUOp_o[0]) );
  AND4X1 U21 ( .A(n13), .B(n5), .C(opcode_i[2]), .D(n12), .Y(Branch_o) );
  CLKBUFX3 U22 ( .A(MemRead_o), .Y(MemToReg_o) );
endmodule


module ALU_DW01_sub_0 ( A, B, CI, DIFF, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] DIFF;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33;
  wire   [32:0] carry;

  XOR3X1 U2_31 ( .A(A[31]), .B(n2), .C(carry[31]), .Y(DIFF[31]) );
  ADDFXL U2_30 ( .A(A[30]), .B(n3), .CI(carry[30]), .CO(carry[31]), .S(
        DIFF[30]) );
  ADDFXL U2_29 ( .A(A[29]), .B(n4), .CI(carry[29]), .CO(carry[30]), .S(
        DIFF[29]) );
  ADDFXL U2_28 ( .A(A[28]), .B(n5), .CI(carry[28]), .CO(carry[29]), .S(
        DIFF[28]) );
  ADDFXL U2_27 ( .A(A[27]), .B(n6), .CI(carry[27]), .CO(carry[28]), .S(
        DIFF[27]) );
  ADDFXL U2_26 ( .A(A[26]), .B(n7), .CI(carry[26]), .CO(carry[27]), .S(
        DIFF[26]) );
  ADDFXL U2_25 ( .A(A[25]), .B(n8), .CI(carry[25]), .CO(carry[26]), .S(
        DIFF[25]) );
  ADDFXL U2_24 ( .A(A[24]), .B(n9), .CI(carry[24]), .CO(carry[25]), .S(
        DIFF[24]) );
  ADDFXL U2_23 ( .A(A[23]), .B(n10), .CI(carry[23]), .CO(carry[24]), .S(
        DIFF[23]) );
  ADDFXL U2_22 ( .A(A[22]), .B(n11), .CI(carry[22]), .CO(carry[23]), .S(
        DIFF[22]) );
  ADDFXL U2_21 ( .A(A[21]), .B(n12), .CI(carry[21]), .CO(carry[22]), .S(
        DIFF[21]) );
  ADDFXL U2_20 ( .A(A[20]), .B(n13), .CI(carry[20]), .CO(carry[21]), .S(
        DIFF[20]) );
  ADDFXL U2_19 ( .A(A[19]), .B(n14), .CI(carry[19]), .CO(carry[20]), .S(
        DIFF[19]) );
  ADDFXL U2_18 ( .A(A[18]), .B(n15), .CI(carry[18]), .CO(carry[19]), .S(
        DIFF[18]) );
  ADDFXL U2_17 ( .A(A[17]), .B(n16), .CI(carry[17]), .CO(carry[18]), .S(
        DIFF[17]) );
  ADDFXL U2_16 ( .A(A[16]), .B(n17), .CI(carry[16]), .CO(carry[17]), .S(
        DIFF[16]) );
  ADDFXL U2_15 ( .A(A[15]), .B(n18), .CI(carry[15]), .CO(carry[16]), .S(
        DIFF[15]) );
  ADDFXL U2_14 ( .A(A[14]), .B(n19), .CI(carry[14]), .CO(carry[15]), .S(
        DIFF[14]) );
  ADDFXL U2_13 ( .A(A[13]), .B(n20), .CI(carry[13]), .CO(carry[14]), .S(
        DIFF[13]) );
  ADDFXL U2_12 ( .A(A[12]), .B(n21), .CI(carry[12]), .CO(carry[13]), .S(
        DIFF[12]) );
  ADDFXL U2_11 ( .A(A[11]), .B(n22), .CI(carry[11]), .CO(carry[12]), .S(
        DIFF[11]) );
  ADDFXL U2_10 ( .A(A[10]), .B(n23), .CI(carry[10]), .CO(carry[11]), .S(
        DIFF[10]) );
  ADDFXL U2_9 ( .A(A[9]), .B(n24), .CI(carry[9]), .CO(carry[10]), .S(DIFF[9])
         );
  ADDFXL U2_8 ( .A(A[8]), .B(n25), .CI(carry[8]), .CO(carry[9]), .S(DIFF[8])
         );
  ADDFXL U2_7 ( .A(A[7]), .B(n26), .CI(carry[7]), .CO(carry[8]), .S(DIFF[7])
         );
  ADDFXL U2_6 ( .A(A[6]), .B(n27), .CI(carry[6]), .CO(carry[7]), .S(DIFF[6])
         );
  ADDFXL U2_5 ( .A(A[5]), .B(n28), .CI(carry[5]), .CO(carry[6]), .S(DIFF[5])
         );
  ADDFXL U2_4 ( .A(A[4]), .B(n29), .CI(carry[4]), .CO(carry[5]), .S(DIFF[4])
         );
  ADDFXL U2_3 ( .A(A[3]), .B(n30), .CI(carry[3]), .CO(carry[4]), .S(DIFF[3])
         );
  ADDFXL U2_2 ( .A(A[2]), .B(n31), .CI(carry[2]), .CO(carry[3]), .S(DIFF[2])
         );
  ADDFXL U2_1 ( .A(A[1]), .B(n32), .CI(carry[1]), .CO(carry[2]), .S(DIFF[1])
         );
  CLKINVX1 U1 ( .A(B[0]), .Y(n33) );
  CLKINVX1 U2 ( .A(B[31]), .Y(n2) );
  NAND2X1 U3 ( .A(B[0]), .B(n1), .Y(carry[1]) );
  CLKINVX1 U4 ( .A(B[1]), .Y(n32) );
  CLKINVX1 U5 ( .A(A[0]), .Y(n1) );
  CLKINVX1 U6 ( .A(B[2]), .Y(n31) );
  CLKINVX1 U7 ( .A(B[3]), .Y(n30) );
  CLKINVX1 U8 ( .A(B[4]), .Y(n29) );
  CLKINVX1 U9 ( .A(B[5]), .Y(n28) );
  CLKINVX1 U10 ( .A(B[6]), .Y(n27) );
  CLKINVX1 U11 ( .A(B[7]), .Y(n26) );
  CLKINVX1 U12 ( .A(B[8]), .Y(n25) );
  CLKINVX1 U13 ( .A(B[9]), .Y(n24) );
  CLKINVX1 U14 ( .A(B[10]), .Y(n23) );
  CLKINVX1 U15 ( .A(B[11]), .Y(n22) );
  CLKINVX1 U16 ( .A(B[12]), .Y(n21) );
  CLKINVX1 U17 ( .A(B[13]), .Y(n20) );
  CLKINVX1 U18 ( .A(B[14]), .Y(n19) );
  CLKINVX1 U19 ( .A(B[15]), .Y(n18) );
  CLKINVX1 U20 ( .A(B[16]), .Y(n17) );
  CLKINVX1 U21 ( .A(B[17]), .Y(n16) );
  CLKINVX1 U22 ( .A(B[18]), .Y(n15) );
  CLKINVX1 U23 ( .A(B[19]), .Y(n14) );
  CLKINVX1 U24 ( .A(B[20]), .Y(n13) );
  CLKINVX1 U25 ( .A(B[21]), .Y(n12) );
  CLKINVX1 U26 ( .A(B[22]), .Y(n11) );
  CLKINVX1 U27 ( .A(B[23]), .Y(n10) );
  CLKINVX1 U28 ( .A(B[24]), .Y(n9) );
  CLKINVX1 U29 ( .A(B[25]), .Y(n8) );
  CLKINVX1 U30 ( .A(B[26]), .Y(n7) );
  CLKINVX1 U31 ( .A(B[27]), .Y(n6) );
  CLKINVX1 U32 ( .A(B[28]), .Y(n5) );
  CLKINVX1 U33 ( .A(B[29]), .Y(n4) );
  CLKINVX1 U34 ( .A(B[30]), .Y(n3) );
  XNOR2X1 U35 ( .A(n33), .B(A[0]), .Y(DIFF[0]) );
endmodule


module ALU_DW01_add_0 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1, n2;
  wire   [31:1] carry;

  ADDFXL U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  ADDFXL U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFXL U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFXL U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFXL U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFXL U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFXL U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFXL U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFXL U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFXL U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFXL U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFXL U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFXL U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFXL U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFXL U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFXL U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFXL U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFXL U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFXL U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFXL U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFXL U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFXL U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  XOR3X1 U1_31 ( .A(A[31]), .B(B[31]), .C(carry[31]), .Y(SUM[31]) );
  ADDFXL U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFXL U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFXL U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXL U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXL U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFXL U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFXL U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFXL U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XNOR2X1 U2 ( .A(B[0]), .B(n2), .Y(SUM[0]) );
  CLKINVX1 U3 ( .A(A[0]), .Y(n2) );
endmodule


module ALU_DW01_cmp6_0 ( A, B, TC, LT, GT, EQ, LE, GE, NE );
  input [31:0] A;
  input [31:0] B;
  input TC;
  output LT, GT, EQ, LE, GE, NE;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104;

  CLKINVX1 U1 ( .A(B[9]), .Y(n22) );
  CLKINVX1 U2 ( .A(B[3]), .Y(n28) );
  CLKINVX1 U3 ( .A(B[2]), .Y(n29) );
  CLKINVX1 U4 ( .A(B[10]), .Y(n21) );
  CLKINVX1 U5 ( .A(B[19]), .Y(n13) );
  CLKINVX1 U6 ( .A(B[21]), .Y(n11) );
  CLKINVX1 U7 ( .A(B[11]), .Y(n20) );
  CLKINVX1 U8 ( .A(B[13]), .Y(n18) );
  CLKINVX1 U9 ( .A(B[20]), .Y(n12) );
  CLKINVX1 U10 ( .A(B[12]), .Y(n19) );
  CLKINVX1 U11 ( .A(B[18]), .Y(n14) );
  CLKINVX1 U12 ( .A(B[26]), .Y(n7) );
  CLKINVX1 U13 ( .A(B[27]), .Y(n5) );
  CLKINVX1 U14 ( .A(B[29]), .Y(n3) );
  CLKINVX1 U15 ( .A(B[28]), .Y(n4) );
  CLKINVX1 U16 ( .A(A[31]), .Y(n1) );
  CLKINVX1 U17 ( .A(B[8]), .Y(n23) );
  CLKINVX1 U18 ( .A(n44), .Y(n6) );
  CLKINVX1 U19 ( .A(n104), .Y(n26) );
  CLKINVX1 U20 ( .A(A[4]), .Y(n27) );
  CLKINVX1 U21 ( .A(A[1]), .Y(n30) );
  CLKINVX1 U22 ( .A(A[7]), .Y(n24) );
  CLKINVX1 U23 ( .A(A[6]), .Y(n25) );
  CLKINVX1 U24 ( .A(A[17]), .Y(n15) );
  CLKINVX1 U25 ( .A(A[16]), .Y(n16) );
  CLKINVX1 U26 ( .A(A[14]), .Y(n17) );
  CLKINVX1 U27 ( .A(B[1]), .Y(n31) );
  CLKINVX1 U28 ( .A(A[25]), .Y(n8) );
  CLKINVX1 U29 ( .A(A[24]), .Y(n9) );
  CLKINVX1 U30 ( .A(A[30]), .Y(n2) );
  CLKINVX1 U31 ( .A(A[22]), .Y(n10) );
  NOR4X1 U32 ( .A(n32), .B(n33), .C(n34), .D(n35), .Y(EQ) );
  NAND4X1 U33 ( .A(n36), .B(n37), .C(n38), .D(n39), .Y(n35) );
  OAI22XL U34 ( .A0(A[1]), .A1(n40), .B0(n40), .B1(n31), .Y(n36) );
  NOR2BX1 U35 ( .AN(A[0]), .B(B[0]), .Y(n40) );
  NAND4BBXL U36 ( .AN(n41), .BN(n42), .C(n43), .D(n44), .Y(n34) );
  NAND2BX1 U37 ( .AN(n45), .B(n46), .Y(n33) );
  NOR4BX1 U38 ( .AN(n47), .B(n48), .C(n49), .D(n50), .Y(n46) );
  NAND4BX1 U39 ( .AN(n51), .B(n52), .C(n53), .D(n54), .Y(n45) );
  NAND4BBXL U40 ( .AN(n55), .BN(n56), .C(n57), .D(n58), .Y(n32) );
  NOR4BBX1 U41 ( .AN(n59), .BN(n60), .C(LT), .D(n61), .Y(n58) );
  OAI22XL U42 ( .A0(B[31]), .A1(n1), .B0(n61), .B1(n62), .Y(LT) );
  AOI32X1 U43 ( .A0(n37), .A1(n38), .A2(n63), .B0(B[30]), .B1(n2), .Y(n62) );
  OAI221XL U44 ( .A0(A[28]), .A1(n4), .B0(A[29]), .B1(n3), .C0(n64), .Y(n63)
         );
  OAI211X1 U45 ( .A0(n65), .A1(n66), .B0(n39), .C0(n43), .Y(n64) );
  NAND2X1 U46 ( .A(A[27]), .B(n5), .Y(n43) );
  NAND2X1 U47 ( .A(A[28]), .B(n4), .Y(n39) );
  OAI32X1 U48 ( .A0(n67), .A1(n41), .A2(n6), .B0(A[26]), .B1(n7), .Y(n66) );
  NAND2X1 U49 ( .A(A[26]), .B(n7), .Y(n44) );
  NOR2X1 U50 ( .A(n8), .B(B[25]), .Y(n41) );
  AOI221XL U51 ( .A0(B[25]), .A1(n8), .B0(B[24]), .B1(n9), .C0(n68), .Y(n67)
         );
  AOI211X1 U52 ( .A0(n69), .A1(n70), .B0(n51), .C0(n42), .Y(n68) );
  NOR2X1 U53 ( .A(n9), .B(B[24]), .Y(n42) );
  NOR2BX1 U54 ( .AN(A[23]), .B(B[23]), .Y(n51) );
  NAND2BX1 U55 ( .AN(A[23]), .B(B[23]), .Y(n70) );
  AOI32X1 U56 ( .A0(n54), .A1(n53), .A2(n71), .B0(B[22]), .B1(n10), .Y(n69) );
  OAI221XL U57 ( .A0(A[20]), .A1(n12), .B0(A[21]), .B1(n11), .C0(n72), .Y(n71)
         );
  OAI211X1 U58 ( .A0(n73), .A1(n74), .B0(n52), .C0(n47), .Y(n72) );
  NAND2X1 U59 ( .A(A[19]), .B(n13), .Y(n47) );
  NAND2X1 U60 ( .A(A[20]), .B(n12), .Y(n52) );
  OAI32X1 U61 ( .A0(n75), .A1(n49), .A2(n50), .B0(A[18]), .B1(n14), .Y(n74) );
  NOR2BX1 U62 ( .AN(A[18]), .B(B[18]), .Y(n50) );
  NOR2X1 U63 ( .A(n15), .B(B[17]), .Y(n49) );
  AOI221XL U64 ( .A0(B[17]), .A1(n15), .B0(B[16]), .B1(n16), .C0(n76), .Y(n75)
         );
  AOI211X1 U65 ( .A0(n77), .A1(n78), .B0(n79), .C0(n48), .Y(n76) );
  NOR2X1 U66 ( .A(n16), .B(B[16]), .Y(n48) );
  NAND2BX1 U67 ( .AN(A[15]), .B(B[15]), .Y(n78) );
  AOI32X1 U68 ( .A0(n80), .A1(n81), .A2(n82), .B0(B[14]), .B1(n17), .Y(n77) );
  OAI221XL U69 ( .A0(A[12]), .A1(n19), .B0(A[13]), .B1(n18), .C0(n83), .Y(n82)
         );
  NAND3X1 U70 ( .A(n84), .B(n85), .C(n86), .Y(n83) );
  OAI221XL U71 ( .A0(A[10]), .A1(n21), .B0(A[11]), .B1(n20), .C0(n87), .Y(n86)
         );
  OAI211X1 U72 ( .A0(n88), .A1(n89), .B0(n90), .C0(n91), .Y(n87) );
  OAI32X1 U73 ( .A0(n92), .A1(n93), .A2(n94), .B0(A[8]), .B1(n23), .Y(n89) );
  AOI221XL U74 ( .A0(B[7]), .A1(n24), .B0(B[6]), .B1(n25), .C0(n95), .Y(n92)
         );
  AOI211X1 U75 ( .A0(n96), .A1(n97), .B0(n98), .C0(n99), .Y(n95) );
  NAND2BX1 U76 ( .AN(A[5]), .B(B[5]), .Y(n97) );
  AOI32X1 U77 ( .A0(n26), .A1(n60), .A2(n100), .B0(B[4]), .B1(n27), .Y(n96) );
  OAI221XL U78 ( .A0(A[2]), .A1(n29), .B0(A[3]), .B1(n28), .C0(n101), .Y(n100)
         );
  OAI211X1 U79 ( .A0(n102), .A1(n30), .B0(n103), .C0(n59), .Y(n101) );
  AO21X1 U80 ( .A0(n30), .A1(n102), .B0(B[1]), .Y(n103) );
  NOR2BX1 U81 ( .AN(B[0]), .B(A[0]), .Y(n102) );
  NOR2X1 U82 ( .A(A[9]), .B(n22), .Y(n88) );
  NOR2X1 U83 ( .A(A[19]), .B(n13), .Y(n73) );
  NAND2X1 U84 ( .A(A[21]), .B(n11), .Y(n53) );
  NAND2BX1 U85 ( .AN(B[22]), .B(A[22]), .Y(n54) );
  NOR2X1 U86 ( .A(A[27]), .B(n5), .Y(n65) );
  OR2X1 U87 ( .A(B[30]), .B(n2), .Y(n38) );
  NAND2X1 U88 ( .A(A[29]), .B(n3), .Y(n37) );
  NOR2BX1 U89 ( .AN(B[31]), .B(A[31]), .Y(n61) );
  NAND2X1 U90 ( .A(A[3]), .B(n28), .Y(n60) );
  NAND2X1 U91 ( .A(A[2]), .B(n29), .Y(n59) );
  NOR4X1 U92 ( .A(n104), .B(n98), .C(n99), .D(n93), .Y(n57) );
  NOR2X1 U93 ( .A(n24), .B(B[7]), .Y(n93) );
  NOR2X1 U94 ( .A(n25), .B(B[6]), .Y(n99) );
  NOR2BX1 U95 ( .AN(A[5]), .B(B[5]), .Y(n98) );
  NOR2X1 U96 ( .A(n27), .B(B[4]), .Y(n104) );
  NAND4BX1 U97 ( .AN(n94), .B(n91), .C(n90), .D(n85), .Y(n56) );
  NAND2X1 U98 ( .A(A[11]), .B(n20), .Y(n85) );
  NAND2X1 U99 ( .A(A[10]), .B(n21), .Y(n90) );
  NAND2X1 U100 ( .A(A[9]), .B(n22), .Y(n91) );
  NOR2BX1 U101 ( .AN(A[8]), .B(B[8]), .Y(n94) );
  NAND4BX1 U102 ( .AN(n79), .B(n84), .C(n81), .D(n80), .Y(n55) );
  NAND2BX1 U103 ( .AN(B[14]), .B(A[14]), .Y(n80) );
  NAND2X1 U104 ( .A(A[13]), .B(n18), .Y(n81) );
  NAND2X1 U105 ( .A(A[12]), .B(n19), .Y(n84) );
  NOR2BX1 U106 ( .AN(A[15]), .B(B[15]), .Y(n79) );
endmodule


module ALU ( ALUCtrl_i, data1_i, data2_i, ALU_o, Zero_o );
  input [3:0] ALUCtrl_i;
  input [31:0] data1_i;
  input [31:0] data2_i;
  output [31:0] ALU_o;
  output Zero_o;
  wire   N107, N108, N109, N110, N111, N112, N113, N114, N115, N116, N117,
         N118, N119, N120, N121, N122, N123, N124, N125, N126, N127, N128,
         N129, N130, N131, N132, N133, N134, N135, N136, N137, N138, N139,
         N140, N141, N142, N143, N144, N145, N146, N147, N148, N149, N150,
         N151, N152, N153, N154, N155, N156, N157, N158, N159, N160, N161,
         N162, N163, N164, N165, N166, N167, N168, N169, N170, N171, n51, n52,
         n53, n54, n55, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107,
         n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118,
         n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129,
         n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140,
         n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151,
         n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162,
         n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173,
         n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n56, n185, n186, n187;

  ALU_DW01_sub_0 sub_371 ( .A(data1_i), .B(data2_i), .CI(1'b0), .DIFF({N170, 
        N169, N168, N167, N166, N165, N164, N163, N162, N161, N160, N159, N158, 
        N157, N156, N155, N154, N153, N152, N151, N150, N149, N148, N147, N146, 
        N145, N144, N143, N142, N141, N140, N139}) );
  ALU_DW01_add_0 add_370 ( .A(data1_i), .B(data2_i), .CI(1'b0), .SUM({N138, 
        N137, N136, N135, N134, N133, N132, N131, N130, N129, N128, N127, N126, 
        N125, N124, N123, N122, N121, N120, N119, N118, N117, N116, N115, N114, 
        N113, N112, N111, N110, N109, N108, N107}) );
  ALU_DW01_cmp6_0 r299 ( .A(data1_i), .B(data2_i), .TC(1'b1), .LT(N171), .EQ(
        Zero_o) );
  CLKINVX1 U5 ( .A(n179), .Y(n185) );
  AND4X1 U6 ( .A(ALUCtrl_i[3]), .B(ALUCtrl_i[2]), .C(n186), .D(n187), .Y(n1)
         );
  CLKBUFX3 U7 ( .A(n58), .Y(n8) );
  CLKBUFX3 U8 ( .A(n58), .Y(n7) );
  CLKBUFX3 U9 ( .A(n185), .Y(n5) );
  CLKBUFX3 U10 ( .A(n185), .Y(n3) );
  CLKBUFX3 U11 ( .A(n185), .Y(n4) );
  CLKBUFX3 U12 ( .A(n58), .Y(n9) );
  CLKBUFX3 U13 ( .A(n185), .Y(n6) );
  OAI211X1 U14 ( .A0(n5), .A1(n44), .B0(n71), .C0(n72), .Y(ALU_o[5]) );
  NAND2X1 U15 ( .A(N112), .B(n7), .Y(n71) );
  AOI221XL U16 ( .A0(N144), .A1(n53), .B0(data2_i[5]), .B1(n73), .C0(n74), .Y(
        n72) );
  OAI21XL U17 ( .A0(n13), .A1(n44), .B0(n4), .Y(n73) );
  OAI211X1 U18 ( .A0(n6), .A1(n41), .B0(n59), .C0(n60), .Y(ALU_o[8]) );
  NAND2X1 U19 ( .A(N115), .B(n7), .Y(n59) );
  AOI221XL U20 ( .A0(N147), .A1(n2), .B0(data2_i[8]), .B1(n61), .C0(n62), .Y(
        n60) );
  OAI21XL U21 ( .A0(n13), .A1(n41), .B0(n5), .Y(n61) );
  OAI21XL U22 ( .A0(n13), .A1(n45), .B0(n5), .Y(n77) );
  OAI21XL U23 ( .A0(n13), .A1(n43), .B0(n5), .Y(n69) );
  OAI21XL U24 ( .A0(n13), .A1(n42), .B0(n5), .Y(n65) );
  OAI211X1 U25 ( .A0(n5), .A1(n47), .B0(n91), .C0(n92), .Y(ALU_o[2]) );
  NAND2X1 U26 ( .A(N109), .B(n7), .Y(n91) );
  AOI221XL U27 ( .A0(N141), .A1(n2), .B0(data2_i[2]), .B1(n93), .C0(n94), .Y(
        n92) );
  OAI21XL U28 ( .A0(n13), .A1(n47), .B0(n4), .Y(n93) );
  OAI211X1 U29 ( .A0(n5), .A1(n46), .B0(n79), .C0(n80), .Y(ALU_o[3]) );
  NAND2X1 U30 ( .A(N110), .B(n7), .Y(n79) );
  AOI221XL U31 ( .A0(N142), .A1(n53), .B0(data2_i[3]), .B1(n81), .C0(n82), .Y(
        n80) );
  OAI21XL U32 ( .A0(n13), .A1(n46), .B0(n5), .Y(n81) );
  CLKINVX1 U33 ( .A(data2_i[0]), .Y(n50) );
  CLKINVX1 U34 ( .A(ALUCtrl_i[2]), .Y(n56) );
  CLKINVX1 U35 ( .A(n1), .Y(n16) );
  CLKINVX1 U36 ( .A(n1), .Y(n17) );
  AND2X2 U37 ( .A(n183), .B(n56), .Y(n58) );
  CLKBUFX3 U38 ( .A(n57), .Y(n14) );
  CLKBUFX3 U39 ( .A(n57), .Y(n13) );
  AND2X2 U40 ( .A(n183), .B(ALUCtrl_i[2]), .Y(n53) );
  AND2X2 U41 ( .A(n183), .B(ALUCtrl_i[2]), .Y(n2) );
  CLKBUFX3 U42 ( .A(n57), .Y(n15) );
  OAI211X1 U43 ( .A0(n5), .A1(n43), .B0(n67), .C0(n68), .Y(ALU_o[6]) );
  NAND2X1 U44 ( .A(N113), .B(n7), .Y(n67) );
  AOI221XL U45 ( .A0(N145), .A1(n2), .B0(data2_i[6]), .B1(n69), .C0(n70), .Y(
        n68) );
  NOR3X1 U46 ( .A(n17), .B(data2_i[6]), .C(data1_i[6]), .Y(n70) );
  OAI211X1 U47 ( .A0(n5), .A1(n42), .B0(n63), .C0(n64), .Y(ALU_o[7]) );
  NAND2X1 U48 ( .A(N114), .B(n7), .Y(n63) );
  AOI221XL U49 ( .A0(N146), .A1(n53), .B0(data2_i[7]), .B1(n65), .C0(n66), .Y(
        n64) );
  NOR3X1 U50 ( .A(n16), .B(data2_i[7]), .C(data1_i[7]), .Y(n66) );
  CLKINVX1 U51 ( .A(data1_i[4]), .Y(n45) );
  CLKINVX1 U52 ( .A(data1_i[6]), .Y(n43) );
  CLKINVX1 U53 ( .A(data1_i[7]), .Y(n42) );
  NOR3X1 U54 ( .A(n17), .B(data2_i[3]), .C(data1_i[3]), .Y(n82) );
  NOR3X1 U55 ( .A(n17), .B(data2_i[2]), .C(data1_i[2]), .Y(n94) );
  NOR3X1 U56 ( .A(n16), .B(data2_i[8]), .C(data1_i[8]), .Y(n62) );
  NOR3X1 U57 ( .A(n17), .B(data2_i[5]), .C(data1_i[5]), .Y(n74) );
  CLKINVX1 U58 ( .A(data1_i[3]), .Y(n46) );
  CLKINVX1 U59 ( .A(data1_i[2]), .Y(n47) );
  CLKINVX1 U60 ( .A(data1_i[8]), .Y(n41) );
  CLKINVX1 U61 ( .A(data1_i[5]), .Y(n44) );
  OAI211X1 U62 ( .A0(n5), .A1(n45), .B0(n75), .C0(n76), .Y(ALU_o[4]) );
  NAND2X1 U63 ( .A(N111), .B(n7), .Y(n75) );
  AOI221XL U64 ( .A0(N143), .A1(n2), .B0(data2_i[4]), .B1(n77), .C0(n78), .Y(
        n76) );
  NOR3X1 U65 ( .A(n16), .B(data2_i[4]), .C(data1_i[4]), .Y(n78) );
  AOI221XL U66 ( .A0(N167), .A1(n2), .B0(data2_i[28]), .B1(n101), .C0(n102), 
        .Y(n100) );
  OAI21XL U67 ( .A0(n13), .A1(n21), .B0(n4), .Y(n101) );
  NOR3X1 U68 ( .A(n17), .B(data2_i[28]), .C(data1_i[28]), .Y(n102) );
  AOI221XL U69 ( .A0(N170), .A1(n2), .B0(data2_i[31]), .B1(n85), .C0(n86), .Y(
        n84) );
  NOR3X1 U70 ( .A(n17), .B(data2_i[31]), .C(data1_i[31]), .Y(n86) );
  OAI21XL U71 ( .A0(n13), .A1(n18), .B0(n4), .Y(n85) );
  AOI221XL U72 ( .A0(N168), .A1(n53), .B0(data2_i[29]), .B1(n97), .C0(n98), 
        .Y(n96) );
  OAI21XL U73 ( .A0(n13), .A1(n20), .B0(n4), .Y(n97) );
  NOR3X1 U74 ( .A(n17), .B(data2_i[29]), .C(data1_i[29]), .Y(n98) );
  AOI221XL U75 ( .A0(N169), .A1(n53), .B0(data2_i[30]), .B1(n89), .C0(n90), 
        .Y(n88) );
  NOR3X1 U76 ( .A(n17), .B(data2_i[30]), .C(data1_i[30]), .Y(n90) );
  OAI21XL U77 ( .A0(n13), .A1(n19), .B0(n5), .Y(n89) );
  AOI33X1 U78 ( .A0(N171), .A1(ALUCtrl_i[1]), .A2(n184), .B0(n49), .B1(n50), 
        .B2(n1), .Y(n181) );
  NOR3X1 U79 ( .A(n186), .B(ALUCtrl_i[3]), .C(n56), .Y(n184) );
  AOI221XL U80 ( .A0(N158), .A1(n2), .B0(data2_i[19]), .B1(n141), .C0(n142), 
        .Y(n140) );
  OAI21XL U81 ( .A0(n14), .A1(n30), .B0(n3), .Y(n141) );
  NOR3X1 U82 ( .A(n16), .B(data2_i[19]), .C(data1_i[19]), .Y(n142) );
  AOI221XL U83 ( .A0(N159), .A1(n2), .B0(data2_i[20]), .B1(n133), .C0(n134), 
        .Y(n132) );
  OAI21XL U84 ( .A0(n14), .A1(n29), .B0(n3), .Y(n133) );
  NOR3X1 U85 ( .A(n16), .B(data2_i[20]), .C(data1_i[20]), .Y(n134) );
  AOI221XL U86 ( .A0(N161), .A1(n2), .B0(data2_i[22]), .B1(n125), .C0(n126), 
        .Y(n124) );
  NOR3X1 U87 ( .A(n17), .B(data2_i[22]), .C(data1_i[22]), .Y(n126) );
  OAI21XL U88 ( .A0(n14), .A1(n27), .B0(n4), .Y(n125) );
  AOI221XL U89 ( .A0(N163), .A1(n2), .B0(data2_i[24]), .B1(n117), .C0(n118), 
        .Y(n116) );
  NOR3X1 U90 ( .A(n17), .B(data2_i[24]), .C(data1_i[24]), .Y(n118) );
  OAI21XL U91 ( .A0(n14), .A1(n25), .B0(n4), .Y(n117) );
  AOI221XL U92 ( .A0(N165), .A1(n2), .B0(data2_i[26]), .B1(n109), .C0(n110), 
        .Y(n108) );
  OAI21XL U93 ( .A0(n14), .A1(n23), .B0(n4), .Y(n109) );
  NOR3X1 U94 ( .A(n17), .B(data2_i[26]), .C(data1_i[26]), .Y(n110) );
  AOI221XL U95 ( .A0(N160), .A1(n53), .B0(data2_i[21]), .B1(n129), .C0(n130), 
        .Y(n128) );
  OAI21XL U96 ( .A0(n14), .A1(n28), .B0(n4), .Y(n129) );
  NOR3X1 U97 ( .A(n17), .B(data2_i[21]), .C(data1_i[21]), .Y(n130) );
  AOI221XL U98 ( .A0(N162), .A1(n53), .B0(data2_i[23]), .B1(n121), .C0(n122), 
        .Y(n120) );
  OAI21XL U99 ( .A0(n14), .A1(n26), .B0(n4), .Y(n121) );
  NOR3X1 U100 ( .A(n17), .B(data2_i[23]), .C(data1_i[23]), .Y(n122) );
  AOI221XL U101 ( .A0(N164), .A1(n53), .B0(data2_i[25]), .B1(n113), .C0(n114), 
        .Y(n112) );
  NOR3X1 U102 ( .A(n17), .B(data2_i[25]), .C(data1_i[25]), .Y(n114) );
  OAI21XL U103 ( .A0(n14), .A1(n24), .B0(n4), .Y(n113) );
  AOI221XL U104 ( .A0(N166), .A1(n53), .B0(data2_i[27]), .B1(n105), .C0(n106), 
        .Y(n104) );
  OAI21XL U105 ( .A0(n13), .A1(n22), .B0(n4), .Y(n105) );
  NOR3X1 U106 ( .A(n17), .B(data2_i[27]), .C(data1_i[27]), .Y(n106) );
  AOI221XL U107 ( .A0(N150), .A1(n2), .B0(data2_i[11]), .B1(n173), .C0(n174), 
        .Y(n172) );
  OAI21XL U108 ( .A0(n15), .A1(n38), .B0(n3), .Y(n173) );
  NOR3X1 U109 ( .A(n16), .B(data2_i[11]), .C(data1_i[11]), .Y(n174) );
  AOI221XL U110 ( .A0(N152), .A1(n2), .B0(data2_i[13]), .B1(n165), .C0(n166), 
        .Y(n164) );
  OAI21XL U111 ( .A0(n15), .A1(n36), .B0(n3), .Y(n165) );
  NOR3X1 U112 ( .A(n16), .B(data2_i[13]), .C(data1_i[13]), .Y(n166) );
  AOI221XL U113 ( .A0(N154), .A1(n2), .B0(data2_i[15]), .B1(n157), .C0(n158), 
        .Y(n156) );
  OAI21XL U114 ( .A0(n14), .A1(n34), .B0(n3), .Y(n157) );
  NOR3X1 U115 ( .A(n16), .B(data2_i[15]), .C(data1_i[15]), .Y(n158) );
  AOI221XL U116 ( .A0(N156), .A1(n2), .B0(data2_i[17]), .B1(n149), .C0(n150), 
        .Y(n148) );
  NOR3X1 U117 ( .A(n16), .B(data2_i[17]), .C(data1_i[17]), .Y(n150) );
  OAI21XL U118 ( .A0(n14), .A1(n32), .B0(n3), .Y(n149) );
  AOI221XL U119 ( .A0(N149), .A1(n53), .B0(data2_i[10]), .B1(n177), .C0(n178), 
        .Y(n176) );
  OAI21XL U120 ( .A0(n15), .A1(n39), .B0(n3), .Y(n177) );
  NOR3X1 U121 ( .A(n16), .B(data2_i[10]), .C(data1_i[10]), .Y(n178) );
  AOI221XL U122 ( .A0(N151), .A1(n53), .B0(data2_i[12]), .B1(n169), .C0(n170), 
        .Y(n168) );
  OAI21XL U123 ( .A0(n15), .A1(n37), .B0(n3), .Y(n169) );
  NOR3X1 U124 ( .A(n16), .B(data2_i[12]), .C(data1_i[12]), .Y(n170) );
  AOI221XL U125 ( .A0(N153), .A1(n53), .B0(data2_i[14]), .B1(n161), .C0(n162), 
        .Y(n160) );
  NOR3X1 U126 ( .A(n16), .B(data2_i[14]), .C(data1_i[14]), .Y(n162) );
  OAI21XL U127 ( .A0(n15), .A1(n35), .B0(n3), .Y(n161) );
  AOI221XL U128 ( .A0(N155), .A1(n53), .B0(data2_i[16]), .B1(n153), .C0(n154), 
        .Y(n152) );
  NOR3X1 U129 ( .A(n16), .B(data2_i[16]), .C(data1_i[16]), .Y(n154) );
  OAI21XL U130 ( .A0(n14), .A1(n33), .B0(n3), .Y(n153) );
  AOI221XL U131 ( .A0(N157), .A1(n53), .B0(data2_i[18]), .B1(n145), .C0(n146), 
        .Y(n144) );
  OAI21XL U132 ( .A0(n14), .A1(n31), .B0(n3), .Y(n145) );
  NOR3X1 U133 ( .A(n16), .B(data2_i[18]), .C(data1_i[18]), .Y(n146) );
  AOI222XL U134 ( .A0(data1_i[0]), .A1(n179), .B0(N139), .B1(n2), .C0(N107), 
        .C1(n9), .Y(n182) );
  AOI221XL U135 ( .A0(N140), .A1(n53), .B0(data2_i[1]), .B1(n137), .C0(n138), 
        .Y(n136) );
  OAI21XL U136 ( .A0(n14), .A1(n48), .B0(n3), .Y(n137) );
  NOR3X1 U137 ( .A(n16), .B(data2_i[1]), .C(data1_i[1]), .Y(n138) );
  AOI221XL U138 ( .A0(N148), .A1(n53), .B0(data2_i[9]), .B1(n54), .C0(n55), 
        .Y(n52) );
  OAI21XL U139 ( .A0(n13), .A1(n40), .B0(n5), .Y(n54) );
  NOR3X1 U140 ( .A(n17), .B(data2_i[9]), .C(data1_i[9]), .Y(n55) );
  CLKINVX1 U141 ( .A(data1_i[14]), .Y(n35) );
  CLKINVX1 U142 ( .A(data1_i[22]), .Y(n27) );
  CLKINVX1 U143 ( .A(data1_i[31]), .Y(n18) );
  CLKINVX1 U144 ( .A(data1_i[1]), .Y(n48) );
  CLKINVX1 U145 ( .A(data1_i[16]), .Y(n33) );
  CLKINVX1 U146 ( .A(data1_i[17]), .Y(n32) );
  CLKINVX1 U147 ( .A(data1_i[24]), .Y(n25) );
  CLKINVX1 U148 ( .A(data1_i[25]), .Y(n24) );
  CLKINVX1 U149 ( .A(data1_i[30]), .Y(n19) );
  CLKINVX1 U150 ( .A(data1_i[9]), .Y(n40) );
  CLKINVX1 U151 ( .A(data1_i[26]), .Y(n23) );
  CLKINVX1 U152 ( .A(data1_i[19]), .Y(n30) );
  CLKINVX1 U153 ( .A(data1_i[27]), .Y(n22) );
  CLKINVX1 U154 ( .A(data1_i[11]), .Y(n38) );
  CLKINVX1 U155 ( .A(data1_i[13]), .Y(n36) );
  CLKINVX1 U156 ( .A(data1_i[21]), .Y(n28) );
  CLKINVX1 U157 ( .A(data1_i[29]), .Y(n20) );
  CLKINVX1 U158 ( .A(data1_i[10]), .Y(n39) );
  CLKINVX1 U159 ( .A(data1_i[12]), .Y(n37) );
  CLKINVX1 U160 ( .A(data1_i[20]), .Y(n29) );
  CLKINVX1 U161 ( .A(data1_i[28]), .Y(n21) );
  CLKINVX1 U162 ( .A(data1_i[18]), .Y(n31) );
  CLKINVX1 U163 ( .A(data1_i[15]), .Y(n34) );
  CLKINVX1 U164 ( .A(data1_i[23]), .Y(n26) );
  CLKINVX1 U165 ( .A(data1_i[0]), .Y(n49) );
  NAND3BX1 U166 ( .AN(ALUCtrl_i[3]), .B(n56), .C(n187), .Y(n57) );
  NOR4X1 U167 ( .A(n186), .B(ALUCtrl_i[1]), .C(ALUCtrl_i[2]), .D(ALUCtrl_i[3]), 
        .Y(n179) );
  NOR3X1 U168 ( .A(ALUCtrl_i[0]), .B(ALUCtrl_i[3]), .C(n187), .Y(n183) );
  CLKINVX1 U169 ( .A(ALUCtrl_i[0]), .Y(n186) );
  CLKINVX1 U170 ( .A(ALUCtrl_i[1]), .Y(n187) );
  OAI211X1 U171 ( .A0(n5), .A1(n48), .B0(n135), .C0(n136), .Y(ALU_o[1]) );
  NAND2X1 U172 ( .A(N108), .B(n8), .Y(n135) );
  OAI211X1 U173 ( .A0(n5), .A1(n34), .B0(n155), .C0(n156), .Y(ALU_o[15]) );
  NAND2X1 U174 ( .A(N122), .B(n8), .Y(n155) );
  OAI211X1 U175 ( .A0(n5), .A1(n33), .B0(n151), .C0(n152), .Y(ALU_o[16]) );
  NAND2X1 U176 ( .A(N123), .B(n8), .Y(n151) );
  OAI211X1 U177 ( .A0(n5), .A1(n32), .B0(n147), .C0(n148), .Y(ALU_o[17]) );
  NAND2X1 U178 ( .A(N124), .B(n8), .Y(n147) );
  OAI211X1 U179 ( .A0(n5), .A1(n31), .B0(n143), .C0(n144), .Y(ALU_o[18]) );
  NAND2X1 U180 ( .A(N125), .B(n8), .Y(n143) );
  OAI211X1 U181 ( .A0(n5), .A1(n30), .B0(n139), .C0(n140), .Y(ALU_o[19]) );
  NAND2X1 U182 ( .A(N126), .B(n8), .Y(n139) );
  OAI211X1 U183 ( .A0(n5), .A1(n29), .B0(n131), .C0(n132), .Y(ALU_o[20]) );
  NAND2X1 U184 ( .A(N127), .B(n8), .Y(n131) );
  OAI211X1 U185 ( .A0(n5), .A1(n28), .B0(n127), .C0(n128), .Y(ALU_o[21]) );
  NAND2X1 U186 ( .A(N128), .B(n8), .Y(n127) );
  OAI211X1 U187 ( .A0(n5), .A1(n27), .B0(n123), .C0(n124), .Y(ALU_o[22]) );
  NAND2X1 U188 ( .A(N129), .B(n8), .Y(n123) );
  OAI211X1 U189 ( .A0(n5), .A1(n26), .B0(n119), .C0(n120), .Y(ALU_o[23]) );
  NAND2X1 U190 ( .A(N130), .B(n8), .Y(n119) );
  OAI211X1 U191 ( .A0(n5), .A1(n25), .B0(n115), .C0(n116), .Y(ALU_o[24]) );
  NAND2X1 U192 ( .A(N131), .B(n8), .Y(n115) );
  OAI211X1 U193 ( .A0(n5), .A1(n24), .B0(n111), .C0(n112), .Y(ALU_o[25]) );
  NAND2X1 U194 ( .A(N132), .B(n8), .Y(n111) );
  OAI211X1 U195 ( .A0(n5), .A1(n23), .B0(n107), .C0(n108), .Y(ALU_o[26]) );
  NAND2X1 U196 ( .A(N133), .B(n8), .Y(n107) );
  OAI211X1 U197 ( .A0(n5), .A1(n22), .B0(n103), .C0(n104), .Y(ALU_o[27]) );
  NAND2X1 U198 ( .A(N134), .B(n7), .Y(n103) );
  OAI211X1 U199 ( .A0(n5), .A1(n21), .B0(n99), .C0(n100), .Y(ALU_o[28]) );
  NAND2X1 U200 ( .A(N135), .B(n7), .Y(n99) );
  OAI211X1 U201 ( .A0(n5), .A1(n20), .B0(n95), .C0(n96), .Y(ALU_o[29]) );
  NAND2X1 U202 ( .A(N136), .B(n7), .Y(n95) );
  OAI211X1 U203 ( .A0(n6), .A1(n39), .B0(n175), .C0(n176), .Y(ALU_o[10]) );
  NAND2X1 U204 ( .A(N117), .B(n9), .Y(n175) );
  OAI211X1 U205 ( .A0(n6), .A1(n38), .B0(n171), .C0(n172), .Y(ALU_o[11]) );
  NAND2X1 U206 ( .A(N118), .B(n9), .Y(n171) );
  OAI211X1 U207 ( .A0(n6), .A1(n37), .B0(n167), .C0(n168), .Y(ALU_o[12]) );
  NAND2X1 U208 ( .A(N119), .B(n9), .Y(n167) );
  OAI211X1 U209 ( .A0(n6), .A1(n36), .B0(n163), .C0(n164), .Y(ALU_o[13]) );
  NAND2X1 U210 ( .A(N120), .B(n9), .Y(n163) );
  OAI211X1 U211 ( .A0(n6), .A1(n35), .B0(n159), .C0(n160), .Y(ALU_o[14]) );
  NAND2X1 U212 ( .A(N121), .B(n9), .Y(n159) );
  OAI211X1 U213 ( .A0(n180), .A1(n50), .B0(n181), .C0(n182), .Y(ALU_o[0]) );
  AOI2BB1X1 U214 ( .A0N(n15), .A1N(n49), .B0(n179), .Y(n180) );
  OAI211X1 U215 ( .A0(n40), .A1(n6), .B0(n51), .C0(n52), .Y(ALU_o[9]) );
  NAND2X1 U216 ( .A(N116), .B(n7), .Y(n51) );
  OAI211X1 U217 ( .A0(n5), .A1(n19), .B0(n87), .C0(n88), .Y(ALU_o[30]) );
  NAND2X1 U218 ( .A(N137), .B(n7), .Y(n87) );
  OAI211X1 U219 ( .A0(n5), .A1(n18), .B0(n83), .C0(n84), .Y(ALU_o[31]) );
  NAND2X1 U220 ( .A(N138), .B(n7), .Y(n83) );
endmodule


module ALUControl ( ALUOp_i, funct_i, ALUctrl_o );
  input [1:0] ALUOp_i;
  input [5:0] funct_i;
  output [3:0] ALUctrl_o;
  wire   n5, n6, n7, n8, n9, n1, n2, n3, n4;

  NOR2X1 U3 ( .A(n5), .B(n1), .Y(ALUctrl_o[3]) );
  CLKINVX1 U4 ( .A(ALUOp_i[1]), .Y(n1) );
  AO22X1 U5 ( .A0(ALUOp_i[0]), .A1(n1), .B0(ALUOp_i[1]), .B1(n6), .Y(
        ALUctrl_o[2]) );
  NAND2X1 U6 ( .A(n7), .B(n3), .Y(n6) );
  AOI222XL U7 ( .A0(funct_i[2]), .A1(funct_i[1]), .B0(funct_i[0]), .B1(n2), 
        .C0(funct_i[3]), .C1(n3), .Y(n5) );
  CLKINVX1 U8 ( .A(funct_i[2]), .Y(n2) );
  AOI21X1 U9 ( .A0(n9), .A1(n7), .B0(n1), .Y(ALUctrl_o[0]) );
  AOI32X1 U10 ( .A0(funct_i[1]), .A1(n4), .A2(funct_i[2]), .B0(funct_i[0]), 
        .B1(n3), .Y(n9) );
  NAND4BX1 U11 ( .AN(funct_i[3]), .B(ALUOp_i[1]), .C(funct_i[2]), .D(n8), .Y(
        ALUctrl_o[1]) );
  NAND2X1 U12 ( .A(funct_i[1]), .B(n4), .Y(n8) );
  AOI2BB1X1 U13 ( .A0N(funct_i[2]), .A1N(n4), .B0(funct_i[3]), .Y(n7) );
  CLKINVX1 U14 ( .A(funct_i[0]), .Y(n4) );
  CLKINVX1 U15 ( .A(funct_i[1]), .Y(n3) );
endmodule


module signExtend ( data_i, data_o );
  input [15:0] data_i;
  output [31:0] data_o;
  wire   data_o_31, n1;
  assign data_o_31 = data_i[15];

  CLKINVX1 U1 ( .A(data_o[25]), .Y(n1) );
  CLKBUFX3 U2 ( .A(data_o_31), .Y(data_o[25]) );
  CLKBUFX3 U3 ( .A(data_o_31), .Y(data_o[30]) );
  CLKBUFX3 U4 ( .A(data_i[14]), .Y(data_o[14]) );
  CLKBUFX3 U5 ( .A(data_i[13]), .Y(data_o[13]) );
  CLKBUFX3 U6 ( .A(data_i[12]), .Y(data_o[12]) );
  CLKBUFX3 U7 ( .A(data_i[11]), .Y(data_o[11]) );
  CLKBUFX3 U8 ( .A(data_i[10]), .Y(data_o[10]) );
  CLKBUFX3 U9 ( .A(data_i[9]), .Y(data_o[9]) );
  CLKBUFX3 U10 ( .A(data_i[8]), .Y(data_o[8]) );
  CLKBUFX3 U11 ( .A(data_i[7]), .Y(data_o[7]) );
  CLKBUFX3 U12 ( .A(data_i[6]), .Y(data_o[6]) );
  CLKBUFX3 U13 ( .A(data_i[5]), .Y(data_o[5]) );
  CLKBUFX3 U14 ( .A(data_i[4]), .Y(data_o[4]) );
  CLKBUFX3 U15 ( .A(data_i[3]), .Y(data_o[3]) );
  CLKBUFX3 U16 ( .A(data_i[2]), .Y(data_o[2]) );
  CLKBUFX3 U17 ( .A(data_i[1]), .Y(data_o[1]) );
  CLKBUFX3 U18 ( .A(data_i[0]), .Y(data_o[0]) );
  CLKINVX1 U19 ( .A(n1), .Y(data_o[29]) );
  CLKINVX1 U20 ( .A(n1), .Y(data_o[28]) );
  CLKINVX1 U21 ( .A(n1), .Y(data_o[27]) );
  CLKINVX1 U22 ( .A(n1), .Y(data_o[31]) );
  CLKINVX1 U23 ( .A(n1), .Y(data_o[24]) );
  CLKINVX1 U24 ( .A(n1), .Y(data_o[23]) );
  CLKINVX1 U25 ( .A(n1), .Y(data_o[22]) );
  CLKINVX1 U26 ( .A(n1), .Y(data_o[21]) );
  CLKINVX1 U27 ( .A(n1), .Y(data_o[20]) );
  CLKINVX1 U28 ( .A(n1), .Y(data_o[19]) );
  CLKINVX1 U29 ( .A(n1), .Y(data_o[18]) );
  CLKINVX1 U30 ( .A(n1), .Y(data_o[17]) );
  CLKINVX1 U31 ( .A(n1), .Y(data_o[16]) );
  CLKINVX1 U32 ( .A(n1), .Y(data_o[15]) );
  CLKINVX1 U33 ( .A(n1), .Y(data_o[26]) );
endmodule


module register_file ( clk, rst, RegWrite_i, WriteReg_i, WriteData_i, 
        ReadReg1_i, ReadReg2_i, ReadData1_o, ReadData2_o, Port28 );
  input [4:0] WriteReg_i;
  input [31:0] WriteData_i;
  input [4:0] ReadReg1_i;
  input [4:0] ReadReg2_i;
  output [31:0] ReadData1_o;
  output [31:0] ReadData2_o;
  input clk, rst, RegWrite_i;
  inout Port28;
  wire   N10, N11, N12, N13, N14, N15, N16, N17, N18, N19, \register[0][31] ,
         \register[0][30] , \register[0][29] , \register[0][28] ,
         \register[0][27] , \register[0][26] , \register[0][25] ,
         \register[0][24] , \register[0][23] , \register[0][22] ,
         \register[0][21] , \register[0][20] , \register[0][19] ,
         \register[0][18] , \register[0][17] , \register[0][16] ,
         \register[0][15] , \register[0][14] , \register[0][13] ,
         \register[0][12] , \register[0][11] , \register[0][10] ,
         \register[0][9] , \register[0][8] , \register[0][7] ,
         \register[0][6] , \register[0][5] , \register[0][4] ,
         \register[0][3] , \register[0][2] , \register[0][1] ,
         \register[0][0] , \register[1][31] , \register[1][30] ,
         \register[1][29] , \register[1][28] , \register[1][27] ,
         \register[1][26] , \register[1][25] , \register[1][24] ,
         \register[1][23] , \register[1][22] , \register[1][21] ,
         \register[1][20] , \register[1][19] , \register[1][18] ,
         \register[1][17] , \register[1][16] , \register[1][15] ,
         \register[1][14] , \register[1][13] , \register[1][12] ,
         \register[1][11] , \register[1][10] , \register[1][9] ,
         \register[1][8] , \register[1][7] , \register[1][6] ,
         \register[1][5] , \register[1][4] , \register[1][3] ,
         \register[1][2] , \register[1][1] , \register[1][0] ,
         \register[2][31] , \register[2][30] , \register[2][29] ,
         \register[2][28] , \register[2][27] , \register[2][26] ,
         \register[2][25] , \register[2][24] , \register[2][23] ,
         \register[2][22] , \register[2][21] , \register[2][20] ,
         \register[2][19] , \register[2][18] , \register[2][17] ,
         \register[2][16] , \register[2][15] , \register[2][14] ,
         \register[2][13] , \register[2][12] , \register[2][11] ,
         \register[2][10] , \register[2][9] , \register[2][8] ,
         \register[2][7] , \register[2][6] , \register[2][5] ,
         \register[2][4] , \register[2][3] , \register[2][2] ,
         \register[2][1] , \register[2][0] , \register[3][31] ,
         \register[3][30] , \register[3][29] , \register[3][28] ,
         \register[3][27] , \register[3][26] , \register[3][25] ,
         \register[3][24] , \register[3][23] , \register[3][22] ,
         \register[3][21] , \register[3][20] , \register[3][19] ,
         \register[3][18] , \register[3][17] , \register[3][16] ,
         \register[3][15] , \register[3][14] , \register[3][13] ,
         \register[3][12] , \register[3][11] , \register[3][10] ,
         \register[3][9] , \register[3][8] , \register[3][7] ,
         \register[3][6] , \register[3][5] , \register[3][4] ,
         \register[3][3] , \register[3][2] , \register[3][1] ,
         \register[3][0] , \register[4][31] , \register[4][30] ,
         \register[4][29] , \register[4][28] , \register[4][27] ,
         \register[4][26] , \register[4][25] , \register[4][24] ,
         \register[4][23] , \register[4][22] , \register[4][21] ,
         \register[4][20] , \register[4][19] , \register[4][18] ,
         \register[4][17] , \register[4][16] , \register[4][15] ,
         \register[4][14] , \register[4][13] , \register[4][12] ,
         \register[4][11] , \register[4][10] , \register[4][9] ,
         \register[4][8] , \register[4][7] , \register[4][6] ,
         \register[4][5] , \register[4][4] , \register[4][3] ,
         \register[4][2] , \register[4][1] , \register[4][0] ,
         \register[5][31] , \register[5][30] , \register[5][29] ,
         \register[5][28] , \register[5][27] , \register[5][26] ,
         \register[5][25] , \register[5][24] , \register[5][23] ,
         \register[5][22] , \register[5][21] , \register[5][20] ,
         \register[5][19] , \register[5][18] , \register[5][17] ,
         \register[5][16] , \register[5][15] , \register[5][14] ,
         \register[5][13] , \register[5][12] , \register[5][11] ,
         \register[5][10] , \register[5][9] , \register[5][8] ,
         \register[5][7] , \register[5][6] , \register[5][5] ,
         \register[5][4] , \register[5][3] , \register[5][2] ,
         \register[5][1] , \register[5][0] , \register[6][31] ,
         \register[6][30] , \register[6][29] , \register[6][28] ,
         \register[6][27] , \register[6][26] , \register[6][25] ,
         \register[6][24] , \register[6][23] , \register[6][22] ,
         \register[6][21] , \register[6][20] , \register[6][19] ,
         \register[6][18] , \register[6][17] , \register[6][16] ,
         \register[6][15] , \register[6][14] , \register[6][13] ,
         \register[6][12] , \register[6][11] , \register[6][10] ,
         \register[6][9] , \register[6][8] , \register[6][7] ,
         \register[6][6] , \register[6][5] , \register[6][4] ,
         \register[6][3] , \register[6][2] , \register[6][1] ,
         \register[6][0] , \register[7][31] , \register[7][30] ,
         \register[7][29] , \register[7][28] , \register[7][27] ,
         \register[7][26] , \register[7][25] , \register[7][24] ,
         \register[7][23] , \register[7][22] , \register[7][21] ,
         \register[7][20] , \register[7][19] , \register[7][18] ,
         \register[7][17] , \register[7][16] , \register[7][15] ,
         \register[7][14] , \register[7][13] , \register[7][12] ,
         \register[7][11] , \register[7][10] , \register[7][9] ,
         \register[7][8] , \register[7][7] , \register[7][6] ,
         \register[7][5] , \register[7][4] , \register[7][3] ,
         \register[7][2] , \register[7][1] , \register[7][0] ,
         \register[8][31] , \register[8][30] , \register[8][29] ,
         \register[8][28] , \register[8][27] , \register[8][26] ,
         \register[8][25] , \register[8][24] , \register[8][23] ,
         \register[8][22] , \register[8][21] , \register[8][20] ,
         \register[8][19] , \register[8][18] , \register[8][17] ,
         \register[8][16] , \register[8][15] , \register[8][14] ,
         \register[8][13] , \register[8][12] , \register[8][11] ,
         \register[8][10] , \register[8][9] , \register[8][8] ,
         \register[8][7] , \register[8][6] , \register[8][5] ,
         \register[8][4] , \register[8][3] , \register[8][2] ,
         \register[8][1] , \register[8][0] , \register[9][31] ,
         \register[9][30] , \register[9][29] , \register[9][28] ,
         \register[9][27] , \register[9][26] , \register[9][25] ,
         \register[9][24] , \register[9][23] , \register[9][22] ,
         \register[9][21] , \register[9][20] , \register[9][19] ,
         \register[9][18] , \register[9][17] , \register[9][16] ,
         \register[9][15] , \register[9][14] , \register[9][13] ,
         \register[9][12] , \register[9][11] , \register[9][10] ,
         \register[9][9] , \register[9][8] , \register[9][7] ,
         \register[9][6] , \register[9][5] , \register[9][4] ,
         \register[9][3] , \register[9][2] , \register[9][1] ,
         \register[9][0] , \register[10][31] , \register[10][30] ,
         \register[10][29] , \register[10][28] , \register[10][27] ,
         \register[10][26] , \register[10][25] , \register[10][24] ,
         \register[10][23] , \register[10][22] , \register[10][21] ,
         \register[10][20] , \register[10][19] , \register[10][18] ,
         \register[10][17] , \register[10][16] , \register[10][15] ,
         \register[10][14] , \register[10][13] , \register[10][12] ,
         \register[10][11] , \register[10][10] , \register[10][9] ,
         \register[10][8] , \register[10][7] , \register[10][6] ,
         \register[10][5] , \register[10][4] , \register[10][3] ,
         \register[10][2] , \register[10][1] , \register[10][0] ,
         \register[11][31] , \register[11][30] , \register[11][29] ,
         \register[11][28] , \register[11][27] , \register[11][26] ,
         \register[11][25] , \register[11][24] , \register[11][23] ,
         \register[11][22] , \register[11][21] , \register[11][20] ,
         \register[11][19] , \register[11][18] , \register[11][17] ,
         \register[11][16] , \register[11][15] , \register[11][14] ,
         \register[11][13] , \register[11][12] , \register[11][11] ,
         \register[11][10] , \register[11][9] , \register[11][8] ,
         \register[11][7] , \register[11][6] , \register[11][5] ,
         \register[11][4] , \register[11][3] , \register[11][2] ,
         \register[11][1] , \register[11][0] , \register[12][31] ,
         \register[12][30] , \register[12][29] , \register[12][28] ,
         \register[12][27] , \register[12][26] , \register[12][25] ,
         \register[12][24] , \register[12][23] , \register[12][22] ,
         \register[12][21] , \register[12][20] , \register[12][19] ,
         \register[12][18] , \register[12][17] , \register[12][16] ,
         \register[12][15] , \register[12][14] , \register[12][13] ,
         \register[12][12] , \register[12][11] , \register[12][10] ,
         \register[12][9] , \register[12][8] , \register[12][7] ,
         \register[12][6] , \register[12][5] , \register[12][4] ,
         \register[12][3] , \register[12][2] , \register[12][1] ,
         \register[12][0] , \register[13][31] , \register[13][30] ,
         \register[13][29] , \register[13][28] , \register[13][27] ,
         \register[13][26] , \register[13][25] , \register[13][24] ,
         \register[13][23] , \register[13][22] , \register[13][21] ,
         \register[13][20] , \register[13][19] , \register[13][18] ,
         \register[13][17] , \register[13][16] , \register[13][15] ,
         \register[13][14] , \register[13][13] , \register[13][12] ,
         \register[13][11] , \register[13][10] , \register[13][9] ,
         \register[13][8] , \register[13][7] , \register[13][6] ,
         \register[13][5] , \register[13][4] , \register[13][3] ,
         \register[13][2] , \register[13][1] , \register[13][0] ,
         \register[14][31] , \register[14][30] , \register[14][29] ,
         \register[14][28] , \register[14][27] , \register[14][26] ,
         \register[14][25] , \register[14][24] , \register[14][23] ,
         \register[14][22] , \register[14][21] , \register[14][20] ,
         \register[14][19] , \register[14][18] , \register[14][17] ,
         \register[14][16] , \register[14][15] , \register[14][14] ,
         \register[14][13] , \register[14][12] , \register[14][11] ,
         \register[14][10] , \register[14][9] , \register[14][8] ,
         \register[14][7] , \register[14][6] , \register[14][5] ,
         \register[14][4] , \register[14][3] , \register[14][2] ,
         \register[14][1] , \register[14][0] , \register[15][31] ,
         \register[15][30] , \register[15][29] , \register[15][28] ,
         \register[15][27] , \register[15][26] , \register[15][25] ,
         \register[15][24] , \register[15][23] , \register[15][22] ,
         \register[15][21] , \register[15][20] , \register[15][19] ,
         \register[15][18] , \register[15][17] , \register[15][16] ,
         \register[15][15] , \register[15][14] , \register[15][13] ,
         \register[15][12] , \register[15][11] , \register[15][10] ,
         \register[15][9] , \register[15][8] , \register[15][7] ,
         \register[15][6] , \register[15][5] , \register[15][4] ,
         \register[15][3] , \register[15][2] , \register[15][1] ,
         \register[15][0] , \register[16][31] , \register[16][30] ,
         \register[16][29] , \register[16][28] , \register[16][27] ,
         \register[16][26] , \register[16][25] , \register[16][24] ,
         \register[16][23] , \register[16][22] , \register[16][21] ,
         \register[16][20] , \register[16][19] , \register[16][18] ,
         \register[16][17] , \register[16][16] , \register[16][15] ,
         \register[16][14] , \register[16][13] , \register[16][12] ,
         \register[16][11] , \register[16][10] , \register[16][9] ,
         \register[16][8] , \register[16][7] , \register[16][6] ,
         \register[16][5] , \register[16][4] , \register[16][3] ,
         \register[16][2] , \register[16][1] , \register[16][0] ,
         \register[17][31] , \register[17][30] , \register[17][29] ,
         \register[17][28] , \register[17][27] , \register[17][26] ,
         \register[17][25] , \register[17][24] , \register[17][23] ,
         \register[17][22] , \register[17][21] , \register[17][20] ,
         \register[17][19] , \register[17][18] , \register[17][17] ,
         \register[17][16] , \register[17][15] , \register[17][14] ,
         \register[17][13] , \register[17][12] , \register[17][11] ,
         \register[17][10] , \register[17][9] , \register[17][8] ,
         \register[17][7] , \register[17][6] , \register[17][5] ,
         \register[17][4] , \register[17][3] , \register[17][2] ,
         \register[17][1] , \register[17][0] , \register[18][31] ,
         \register[18][30] , \register[18][29] , \register[18][28] ,
         \register[18][27] , \register[18][26] , \register[18][25] ,
         \register[18][24] , \register[18][23] , \register[18][22] ,
         \register[18][21] , \register[18][20] , \register[18][19] ,
         \register[18][18] , \register[18][17] , \register[18][16] ,
         \register[18][15] , \register[18][14] , \register[18][13] ,
         \register[18][12] , \register[18][11] , \register[18][10] ,
         \register[18][9] , \register[18][8] , \register[18][7] ,
         \register[18][6] , \register[18][5] , \register[18][4] ,
         \register[18][3] , \register[18][2] , \register[18][1] ,
         \register[18][0] , \register[19][31] , \register[19][30] ,
         \register[19][29] , \register[19][28] , \register[19][27] ,
         \register[19][26] , \register[19][25] , \register[19][24] ,
         \register[19][23] , \register[19][22] , \register[19][21] ,
         \register[19][20] , \register[19][19] , \register[19][18] ,
         \register[19][17] , \register[19][16] , \register[19][15] ,
         \register[19][14] , \register[19][13] , \register[19][12] ,
         \register[19][11] , \register[19][10] , \register[19][9] ,
         \register[19][8] , \register[19][7] , \register[19][6] ,
         \register[19][5] , \register[19][4] , \register[19][3] ,
         \register[19][2] , \register[19][1] , \register[19][0] ,
         \register[20][31] , \register[20][30] , \register[20][29] ,
         \register[20][28] , \register[20][27] , \register[20][26] ,
         \register[20][25] , \register[20][24] , \register[20][23] ,
         \register[20][22] , \register[20][21] , \register[20][20] ,
         \register[20][19] , \register[20][18] , \register[20][17] ,
         \register[20][16] , \register[20][15] , \register[20][14] ,
         \register[20][13] , \register[20][12] , \register[20][11] ,
         \register[20][10] , \register[20][9] , \register[20][8] ,
         \register[20][7] , \register[20][6] , \register[20][5] ,
         \register[20][4] , \register[20][3] , \register[20][2] ,
         \register[20][1] , \register[20][0] , \register[21][31] ,
         \register[21][30] , \register[21][29] , \register[21][28] ,
         \register[21][27] , \register[21][26] , \register[21][25] ,
         \register[21][24] , \register[21][23] , \register[21][22] ,
         \register[21][21] , \register[21][20] , \register[21][19] ,
         \register[21][18] , \register[21][17] , \register[21][16] ,
         \register[21][15] , \register[21][14] , \register[21][13] ,
         \register[21][12] , \register[21][11] , \register[21][10] ,
         \register[21][9] , \register[21][8] , \register[21][7] ,
         \register[21][6] , \register[21][5] , \register[21][4] ,
         \register[21][3] , \register[21][2] , \register[21][1] ,
         \register[21][0] , \register[22][31] , \register[22][30] ,
         \register[22][29] , \register[22][28] , \register[22][27] ,
         \register[22][26] , \register[22][25] , \register[22][24] ,
         \register[22][23] , \register[22][22] , \register[22][21] ,
         \register[22][20] , \register[22][19] , \register[22][18] ,
         \register[22][17] , \register[22][16] , \register[22][15] ,
         \register[22][14] , \register[22][13] , \register[22][12] ,
         \register[22][11] , \register[22][10] , \register[22][9] ,
         \register[22][8] , \register[22][7] , \register[22][6] ,
         \register[22][5] , \register[22][4] , \register[22][3] ,
         \register[22][2] , \register[22][1] , \register[22][0] ,
         \register[23][31] , \register[23][30] , \register[23][29] ,
         \register[23][28] , \register[23][27] , \register[23][26] ,
         \register[23][25] , \register[23][24] , \register[23][23] ,
         \register[23][22] , \register[23][21] , \register[23][20] ,
         \register[23][19] , \register[23][18] , \register[23][17] ,
         \register[23][16] , \register[23][15] , \register[23][14] ,
         \register[23][13] , \register[23][12] , \register[23][11] ,
         \register[23][10] , \register[23][9] , \register[23][8] ,
         \register[23][7] , \register[23][6] , \register[23][5] ,
         \register[23][4] , \register[23][3] , \register[23][2] ,
         \register[23][1] , \register[23][0] , \register[24][31] ,
         \register[24][30] , \register[24][29] , \register[24][28] ,
         \register[24][27] , \register[24][26] , \register[24][25] ,
         \register[24][24] , \register[24][23] , \register[24][22] ,
         \register[24][21] , \register[24][20] , \register[24][19] ,
         \register[24][18] , \register[24][17] , \register[24][16] ,
         \register[24][15] , \register[24][14] , \register[24][13] ,
         \register[24][12] , \register[24][11] , \register[24][10] ,
         \register[24][9] , \register[24][8] , \register[24][7] ,
         \register[24][6] , \register[24][5] , \register[24][4] ,
         \register[24][3] , \register[24][2] , \register[24][1] ,
         \register[24][0] , \register[25][31] , \register[25][30] ,
         \register[25][29] , \register[25][28] , \register[25][27] ,
         \register[25][26] , \register[25][25] , \register[25][24] ,
         \register[25][23] , \register[25][22] , \register[25][21] ,
         \register[25][20] , \register[25][19] , \register[25][18] ,
         \register[25][17] , \register[25][16] , \register[25][15] ,
         \register[25][14] , \register[25][13] , \register[25][12] ,
         \register[25][11] , \register[25][10] , \register[25][9] ,
         \register[25][8] , \register[25][7] , \register[25][6] ,
         \register[25][5] , \register[25][4] , \register[25][3] ,
         \register[25][2] , \register[25][1] , \register[25][0] ,
         \register[26][31] , \register[26][30] , \register[26][29] ,
         \register[26][28] , \register[26][27] , \register[26][26] ,
         \register[26][25] , \register[26][24] , \register[26][23] ,
         \register[26][22] , \register[26][21] , \register[26][20] ,
         \register[26][19] , \register[26][18] , \register[26][17] ,
         \register[26][16] , \register[26][15] , \register[26][14] ,
         \register[26][13] , \register[26][12] , \register[26][11] ,
         \register[26][10] , \register[26][9] , \register[26][8] ,
         \register[26][7] , \register[26][6] , \register[26][5] ,
         \register[26][4] , \register[26][3] , \register[26][2] ,
         \register[26][1] , \register[26][0] , \register[27][31] ,
         \register[27][30] , \register[27][29] , \register[27][28] ,
         \register[27][27] , \register[27][26] , \register[27][25] ,
         \register[27][24] , \register[27][23] , \register[27][22] ,
         \register[27][21] , \register[27][20] , \register[27][19] ,
         \register[27][18] , \register[27][17] , \register[27][16] ,
         \register[27][15] , \register[27][14] , \register[27][13] ,
         \register[27][12] , \register[27][11] , \register[27][10] ,
         \register[27][9] , \register[27][8] , \register[27][7] ,
         \register[27][6] , \register[27][5] , \register[27][4] ,
         \register[27][3] , \register[27][2] , \register[27][1] ,
         \register[27][0] , \register[28][31] , \register[28][30] ,
         \register[28][29] , \register[28][28] , \register[28][27] ,
         \register[28][26] , \register[28][25] , \register[28][24] ,
         \register[28][23] , \register[28][22] , \register[28][21] ,
         \register[28][20] , \register[28][19] , \register[28][18] ,
         \register[28][17] , \register[28][16] , \register[28][15] ,
         \register[28][14] , \register[28][13] , \register[28][12] ,
         \register[28][11] , \register[28][10] , \register[28][9] ,
         \register[28][8] , \register[28][7] , \register[28][6] ,
         \register[28][5] , \register[28][4] , \register[28][3] ,
         \register[28][2] , \register[28][1] , \register[28][0] ,
         \register[29][31] , \register[29][30] , \register[29][29] ,
         \register[29][28] , \register[29][27] , \register[29][26] ,
         \register[29][25] , \register[29][24] , \register[29][23] ,
         \register[29][22] , \register[29][21] , \register[29][20] ,
         \register[29][19] , \register[29][18] , \register[29][17] ,
         \register[29][16] , \register[29][15] , \register[29][14] ,
         \register[29][13] , \register[29][12] , \register[29][11] ,
         \register[29][10] , \register[29][9] , \register[29][8] ,
         \register[29][7] , \register[29][6] , \register[29][5] ,
         \register[29][4] , \register[29][3] , \register[29][2] ,
         \register[29][1] , \register[29][0] , \register[30][31] ,
         \register[30][30] , \register[30][29] , \register[30][28] ,
         \register[30][27] , \register[30][26] , \register[30][25] ,
         \register[30][24] , \register[30][23] , \register[30][22] ,
         \register[30][21] , \register[30][20] , \register[30][19] ,
         \register[30][18] , \register[30][17] , \register[30][16] ,
         \register[30][15] , \register[30][14] , \register[30][13] ,
         \register[30][12] , \register[30][11] , \register[30][10] ,
         \register[30][9] , \register[30][8] , \register[30][7] ,
         \register[30][6] , \register[30][5] , \register[30][4] ,
         \register[30][3] , \register[30][2] , \register[30][1] ,
         \register[30][0] , \register[31][31] , \register[31][30] ,
         \register[31][29] , \register[31][28] , \register[31][27] ,
         \register[31][26] , \register[31][25] , \register[31][24] ,
         \register[31][23] , \register[31][22] , \register[31][21] ,
         \register[31][20] , \register[31][19] , \register[31][18] ,
         \register[31][17] , \register[31][16] , \register[31][15] ,
         \register[31][14] , \register[31][13] , \register[31][12] ,
         \register[31][11] , \register[31][10] , \register[31][9] ,
         \register[31][8] , \register[31][7] , \register[31][6] ,
         \register[31][5] , \register[31][4] , \register[31][3] ,
         \register[31][2] , \register[31][1] , \register[31][0] , n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107,
         n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118,
         n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129,
         n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140,
         n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151,
         n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162,
         n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173,
         n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184,
         n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195,
         n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206,
         n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217,
         n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228,
         n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239,
         n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250,
         n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261,
         n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272,
         n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283,
         n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294,
         n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
         n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316,
         n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327,
         n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338,
         n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349,
         n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
         n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
         n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
         n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
         n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
         n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
         n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
         n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
         n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
         n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
         n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
         n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
         n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
         n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038,
         n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048,
         n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058,
         n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068,
         n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078,
         n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
         n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
         n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1, n2, n3, n4, n5,
         n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
         n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
         n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
         n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
         n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
         n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
         n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
         n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
         n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
         n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
         n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
         n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
         n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
         n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
         n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
         n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
         n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
         n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
         n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
         n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303,
         n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313,
         n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323,
         n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333,
         n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343,
         n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353,
         n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363,
         n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373,
         n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383,
         n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393,
         n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403,
         n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413,
         n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423,
         n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433,
         n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443,
         n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453,
         n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463,
         n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473,
         n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483,
         n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493,
         n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503,
         n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513,
         n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523,
         n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533,
         n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543,
         n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553,
         n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563,
         n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573,
         n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583,
         n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593,
         n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603,
         n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613,
         n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623,
         n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633,
         n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643,
         n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653,
         n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663,
         n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673,
         n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683,
         n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693,
         n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703,
         n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713,
         n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723,
         n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733,
         n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743,
         n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753,
         n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763,
         n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773,
         n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783,
         n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793,
         n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803,
         n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813,
         n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823,
         n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833,
         n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843,
         n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853,
         n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863,
         n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873,
         n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883,
         n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893,
         n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903,
         n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913,
         n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923,
         n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933,
         n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943,
         n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953,
         n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963,
         n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973,
         n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983,
         n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993,
         n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003,
         n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013,
         n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023,
         n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033,
         n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043,
         n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053,
         n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063,
         n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073,
         n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083,
         n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093,
         n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103,
         n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113,
         n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123,
         n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133,
         n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143,
         n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153,
         n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163,
         n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173,
         n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183,
         n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193,
         n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203,
         n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213,
         n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223,
         n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233,
         n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243,
         n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253,
         n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263,
         n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273,
         n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283,
         n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293,
         n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303,
         n2304, n2305, n2306, n2307, n2308, n2309, n2310;
  assign N10 = ReadReg1_i[0];
  assign N11 = ReadReg1_i[1];
  assign N12 = ReadReg1_i[2];
  assign N13 = ReadReg1_i[3];
  assign N14 = ReadReg1_i[4];
  assign N15 = ReadReg2_i[0];
  assign N16 = ReadReg2_i[1];
  assign N17 = ReadReg2_i[2];
  assign N18 = ReadReg2_i[3];
  assign N19 = ReadReg2_i[4];

  DFFRX1 \register_reg[3][31]  ( .D(n1009), .CK(clk), .RN(n2098), .Q(
        \register[3][31] ) );
  DFFRX1 \register_reg[3][30]  ( .D(n1008), .CK(clk), .RN(n2098), .Q(
        \register[3][30] ) );
  DFFRX1 \register_reg[3][29]  ( .D(n1007), .CK(clk), .RN(n2098), .Q(
        \register[3][29] ) );
  DFFRX1 \register_reg[3][28]  ( .D(n1006), .CK(clk), .RN(n2098), .Q(
        \register[3][28] ) );
  DFFRX1 \register_reg[3][27]  ( .D(n1005), .CK(clk), .RN(n2098), .Q(
        \register[3][27] ) );
  DFFRX1 \register_reg[3][26]  ( .D(n1004), .CK(clk), .RN(n2097), .Q(
        \register[3][26] ) );
  DFFRX1 \register_reg[3][25]  ( .D(n1003), .CK(clk), .RN(n2097), .Q(
        \register[3][25] ) );
  DFFRX1 \register_reg[3][24]  ( .D(n1002), .CK(clk), .RN(n2097), .Q(
        \register[3][24] ) );
  DFFRX1 \register_reg[3][23]  ( .D(n1001), .CK(clk), .RN(n2097), .Q(
        \register[3][23] ) );
  DFFRX1 \register_reg[3][22]  ( .D(n1000), .CK(clk), .RN(n2097), .Q(
        \register[3][22] ) );
  DFFRX1 \register_reg[3][21]  ( .D(n999), .CK(clk), .RN(n2097), .Q(
        \register[3][21] ) );
  DFFRX1 \register_reg[3][20]  ( .D(n998), .CK(clk), .RN(n2097), .Q(
        \register[3][20] ) );
  DFFRX1 \register_reg[3][19]  ( .D(n997), .CK(clk), .RN(n2097), .Q(
        \register[3][19] ) );
  DFFRX1 \register_reg[3][18]  ( .D(n996), .CK(clk), .RN(n2097), .Q(
        \register[3][18] ) );
  DFFRX1 \register_reg[3][17]  ( .D(n995), .CK(clk), .RN(n2097), .Q(
        \register[3][17] ) );
  DFFRX1 \register_reg[3][16]  ( .D(n994), .CK(clk), .RN(n2097), .Q(
        \register[3][16] ) );
  DFFRX1 \register_reg[3][15]  ( .D(n993), .CK(clk), .RN(n2097), .Q(
        \register[3][15] ) );
  DFFRX1 \register_reg[3][14]  ( .D(n992), .CK(clk), .RN(n2097), .Q(
        \register[3][14] ) );
  DFFRX1 \register_reg[3][13]  ( .D(n991), .CK(clk), .RN(n2096), .Q(
        \register[3][13] ) );
  DFFRX1 \register_reg[3][12]  ( .D(n990), .CK(clk), .RN(n2096), .Q(
        \register[3][12] ) );
  DFFRX1 \register_reg[3][11]  ( .D(n989), .CK(clk), .RN(n2096), .Q(
        \register[3][11] ) );
  DFFRX1 \register_reg[3][10]  ( .D(n988), .CK(clk), .RN(n2096), .Q(
        \register[3][10] ) );
  DFFRX1 \register_reg[3][9]  ( .D(n987), .CK(clk), .RN(n2096), .Q(
        \register[3][9] ) );
  DFFRX1 \register_reg[7][31]  ( .D(n881), .CK(clk), .RN(n2088), .Q(
        \register[7][31] ) );
  DFFRX1 \register_reg[7][30]  ( .D(n880), .CK(clk), .RN(n2088), .Q(
        \register[7][30] ) );
  DFFRX1 \register_reg[7][29]  ( .D(n879), .CK(clk), .RN(n2088), .Q(
        \register[7][29] ) );
  DFFRX1 \register_reg[7][28]  ( .D(n878), .CK(clk), .RN(n2088), .Q(
        \register[7][28] ) );
  DFFRX1 \register_reg[7][27]  ( .D(n877), .CK(clk), .RN(n2088), .Q(
        \register[7][27] ) );
  DFFRX1 \register_reg[7][26]  ( .D(n876), .CK(clk), .RN(n2088), .Q(
        \register[7][26] ) );
  DFFRX1 \register_reg[7][25]  ( .D(n875), .CK(clk), .RN(n2088), .Q(
        \register[7][25] ) );
  DFFRX1 \register_reg[7][24]  ( .D(n874), .CK(clk), .RN(n2087), .Q(
        \register[7][24] ) );
  DFFRX1 \register_reg[7][23]  ( .D(n873), .CK(clk), .RN(n2087), .Q(
        \register[7][23] ) );
  DFFRX1 \register_reg[7][22]  ( .D(n872), .CK(clk), .RN(n2087), .Q(
        \register[7][22] ) );
  DFFRX1 \register_reg[7][21]  ( .D(n871), .CK(clk), .RN(n2087), .Q(
        \register[7][21] ) );
  DFFRX1 \register_reg[7][20]  ( .D(n870), .CK(clk), .RN(n2087), .Q(
        \register[7][20] ) );
  DFFRX1 \register_reg[7][19]  ( .D(n869), .CK(clk), .RN(n2087), .Q(
        \register[7][19] ) );
  DFFRX1 \register_reg[7][18]  ( .D(n868), .CK(clk), .RN(n2087), .Q(
        \register[7][18] ) );
  DFFRX1 \register_reg[7][17]  ( .D(n867), .CK(clk), .RN(n2087), .Q(
        \register[7][17] ) );
  DFFRX1 \register_reg[7][16]  ( .D(n866), .CK(clk), .RN(n2087), .Q(
        \register[7][16] ) );
  DFFRX1 \register_reg[7][15]  ( .D(n865), .CK(clk), .RN(n2087), .Q(
        \register[7][15] ) );
  DFFRX1 \register_reg[7][14]  ( .D(n864), .CK(clk), .RN(n2087), .Q(
        \register[7][14] ) );
  DFFRX1 \register_reg[7][13]  ( .D(n863), .CK(clk), .RN(n2087), .Q(
        \register[7][13] ) );
  DFFRX1 \register_reg[7][12]  ( .D(n862), .CK(clk), .RN(n2087), .Q(
        \register[7][12] ) );
  DFFRX1 \register_reg[7][11]  ( .D(n861), .CK(clk), .RN(n2086), .Q(
        \register[7][11] ) );
  DFFRX1 \register_reg[7][10]  ( .D(n860), .CK(clk), .RN(n2086), .Q(
        \register[7][10] ) );
  DFFRX1 \register_reg[7][9]  ( .D(n859), .CK(clk), .RN(n2086), .Q(
        \register[7][9] ) );
  DFFRX1 \register_reg[11][31]  ( .D(n753), .CK(clk), .RN(n2078), .Q(
        \register[11][31] ) );
  DFFRX1 \register_reg[11][30]  ( .D(n752), .CK(clk), .RN(n2078), .Q(
        \register[11][30] ) );
  DFFRX1 \register_reg[11][29]  ( .D(n751), .CK(clk), .RN(n2078), .Q(
        \register[11][29] ) );
  DFFRX1 \register_reg[11][28]  ( .D(n750), .CK(clk), .RN(n2078), .Q(
        \register[11][28] ) );
  DFFRX1 \register_reg[11][27]  ( .D(n749), .CK(clk), .RN(n2078), .Q(
        \register[11][27] ) );
  DFFRX1 \register_reg[11][26]  ( .D(n748), .CK(clk), .RN(n2078), .Q(
        \register[11][26] ) );
  DFFRX1 \register_reg[11][25]  ( .D(n747), .CK(clk), .RN(n2078), .Q(
        \register[11][25] ) );
  DFFRX1 \register_reg[11][24]  ( .D(n746), .CK(clk), .RN(n2078), .Q(
        \register[11][24] ) );
  DFFRX1 \register_reg[11][23]  ( .D(n745), .CK(clk), .RN(n2078), .Q(
        \register[11][23] ) );
  DFFRX1 \register_reg[11][22]  ( .D(n744), .CK(clk), .RN(n2077), .Q(
        \register[11][22] ) );
  DFFRX1 \register_reg[11][21]  ( .D(n743), .CK(clk), .RN(n2077), .Q(
        \register[11][21] ) );
  DFFRX1 \register_reg[11][20]  ( .D(n742), .CK(clk), .RN(n2077), .Q(
        \register[11][20] ) );
  DFFRX1 \register_reg[11][19]  ( .D(n741), .CK(clk), .RN(n2077), .Q(
        \register[11][19] ) );
  DFFRX1 \register_reg[11][18]  ( .D(n740), .CK(clk), .RN(n2077), .Q(
        \register[11][18] ) );
  DFFRX1 \register_reg[11][17]  ( .D(n739), .CK(clk), .RN(n2077), .Q(
        \register[11][17] ) );
  DFFRX1 \register_reg[11][16]  ( .D(n738), .CK(clk), .RN(n2077), .Q(
        \register[11][16] ) );
  DFFRX1 \register_reg[11][15]  ( .D(n737), .CK(clk), .RN(n2077), .Q(
        \register[11][15] ) );
  DFFRX1 \register_reg[11][14]  ( .D(n736), .CK(clk), .RN(n2077), .Q(
        \register[11][14] ) );
  DFFRX1 \register_reg[11][13]  ( .D(n735), .CK(clk), .RN(n2077), .Q(
        \register[11][13] ) );
  DFFRX1 \register_reg[11][12]  ( .D(n734), .CK(clk), .RN(n2077), .Q(
        \register[11][12] ) );
  DFFRX1 \register_reg[11][11]  ( .D(n733), .CK(clk), .RN(n2077), .Q(
        \register[11][11] ) );
  DFFRX1 \register_reg[11][10]  ( .D(n732), .CK(clk), .RN(n2077), .Q(
        \register[11][10] ) );
  DFFRX1 \register_reg[11][9]  ( .D(n731), .CK(clk), .RN(n2076), .Q(
        \register[11][9] ) );
  DFFRX1 \register_reg[15][31]  ( .D(n625), .CK(clk), .RN(n2068), .Q(
        \register[15][31] ) );
  DFFRX1 \register_reg[15][30]  ( .D(n624), .CK(clk), .RN(n2068), .Q(
        \register[15][30] ) );
  DFFRX1 \register_reg[15][29]  ( .D(n623), .CK(clk), .RN(n2068), .Q(
        \register[15][29] ) );
  DFFRX1 \register_reg[15][28]  ( .D(n622), .CK(clk), .RN(n2068), .Q(
        \register[15][28] ) );
  DFFRX1 \register_reg[15][27]  ( .D(n621), .CK(clk), .RN(n2068), .Q(
        \register[15][27] ) );
  DFFRX1 \register_reg[15][26]  ( .D(n620), .CK(clk), .RN(n2068), .Q(
        \register[15][26] ) );
  DFFRX1 \register_reg[15][25]  ( .D(n619), .CK(clk), .RN(n2068), .Q(
        \register[15][25] ) );
  DFFRX1 \register_reg[15][24]  ( .D(n618), .CK(clk), .RN(n2068), .Q(
        \register[15][24] ) );
  DFFRX1 \register_reg[15][23]  ( .D(n617), .CK(clk), .RN(n2068), .Q(
        \register[15][23] ) );
  DFFRX1 \register_reg[15][22]  ( .D(n616), .CK(clk), .RN(n2068), .Q(
        \register[15][22] ) );
  DFFRX1 \register_reg[15][21]  ( .D(n615), .CK(clk), .RN(n2068), .Q(
        \register[15][21] ) );
  DFFRX1 \register_reg[15][20]  ( .D(n614), .CK(clk), .RN(n2067), .Q(
        \register[15][20] ) );
  DFFRX1 \register_reg[15][19]  ( .D(n613), .CK(clk), .RN(n2067), .Q(
        \register[15][19] ) );
  DFFRX1 \register_reg[15][18]  ( .D(n612), .CK(clk), .RN(n2067), .Q(
        \register[15][18] ) );
  DFFRX1 \register_reg[15][17]  ( .D(n611), .CK(clk), .RN(n2067), .Q(
        \register[15][17] ) );
  DFFRX1 \register_reg[15][16]  ( .D(n610), .CK(clk), .RN(n2067), .Q(
        \register[15][16] ) );
  DFFRX1 \register_reg[15][15]  ( .D(n609), .CK(clk), .RN(n2067), .Q(
        \register[15][15] ) );
  DFFRX1 \register_reg[15][14]  ( .D(n608), .CK(clk), .RN(n2067), .Q(
        \register[15][14] ) );
  DFFRX1 \register_reg[15][13]  ( .D(n607), .CK(clk), .RN(n2067), .Q(
        \register[15][13] ) );
  DFFRX1 \register_reg[15][12]  ( .D(n606), .CK(clk), .RN(n2067), .Q(
        \register[15][12] ) );
  DFFRX1 \register_reg[15][11]  ( .D(n605), .CK(clk), .RN(n2067), .Q(
        \register[15][11] ) );
  DFFRX1 \register_reg[15][10]  ( .D(n604), .CK(clk), .RN(n2067), .Q(
        \register[15][10] ) );
  DFFRX1 \register_reg[15][9]  ( .D(n603), .CK(clk), .RN(n2067), .Q(
        \register[15][9] ) );
  DFFRX1 \register_reg[19][31]  ( .D(n497), .CK(clk), .RN(n2058), .Q(
        \register[19][31] ) );
  DFFRX1 \register_reg[19][30]  ( .D(n496), .CK(clk), .RN(n2058), .Q(
        \register[19][30] ) );
  DFFRX1 \register_reg[19][29]  ( .D(n495), .CK(clk), .RN(n2058), .Q(
        \register[19][29] ) );
  DFFRX1 \register_reg[19][28]  ( .D(n494), .CK(clk), .RN(n2058), .Q(
        \register[19][28] ) );
  DFFRX1 \register_reg[19][27]  ( .D(n493), .CK(clk), .RN(n2058), .Q(
        \register[19][27] ) );
  DFFRX1 \register_reg[19][26]  ( .D(n492), .CK(clk), .RN(n2058), .Q(
        \register[19][26] ) );
  DFFRX1 \register_reg[19][25]  ( .D(n491), .CK(clk), .RN(n2058), .Q(
        \register[19][25] ) );
  DFFRX1 \register_reg[19][24]  ( .D(n490), .CK(clk), .RN(n2058), .Q(
        \register[19][24] ) );
  DFFRX1 \register_reg[19][23]  ( .D(n489), .CK(clk), .RN(n2058), .Q(
        \register[19][23] ) );
  DFFRX1 \register_reg[19][22]  ( .D(n488), .CK(clk), .RN(n2058), .Q(
        \register[19][22] ) );
  DFFRX1 \register_reg[19][21]  ( .D(n487), .CK(clk), .RN(n2058), .Q(
        \register[19][21] ) );
  DFFRX1 \register_reg[19][20]  ( .D(n486), .CK(clk), .RN(n2058), .Q(
        \register[19][20] ) );
  DFFRX1 \register_reg[19][19]  ( .D(n485), .CK(clk), .RN(n2058), .Q(
        \register[19][19] ) );
  DFFRX1 \register_reg[19][18]  ( .D(n484), .CK(clk), .RN(n2057), .Q(
        \register[19][18] ) );
  DFFRX1 \register_reg[19][17]  ( .D(n483), .CK(clk), .RN(n2057), .Q(
        \register[19][17] ) );
  DFFRX1 \register_reg[19][16]  ( .D(n482), .CK(clk), .RN(n2057), .Q(
        \register[19][16] ) );
  DFFRX1 \register_reg[19][15]  ( .D(n481), .CK(clk), .RN(n2057), .Q(
        \register[19][15] ) );
  DFFRX1 \register_reg[19][14]  ( .D(n480), .CK(clk), .RN(n2057), .Q(
        \register[19][14] ) );
  DFFRX1 \register_reg[19][13]  ( .D(n479), .CK(clk), .RN(n2057), .Q(
        \register[19][13] ) );
  DFFRX1 \register_reg[19][12]  ( .D(n478), .CK(clk), .RN(n2057), .Q(
        \register[19][12] ) );
  DFFRX1 \register_reg[19][11]  ( .D(n477), .CK(clk), .RN(n2057), .Q(
        \register[19][11] ) );
  DFFRX1 \register_reg[19][10]  ( .D(n476), .CK(clk), .RN(n2057), .Q(
        \register[19][10] ) );
  DFFRX1 \register_reg[19][9]  ( .D(n475), .CK(clk), .RN(n2057), .Q(
        \register[19][9] ) );
  DFFRX1 \register_reg[23][31]  ( .D(n369), .CK(clk), .RN(n2049), .Q(
        \register[23][31] ) );
  DFFRX1 \register_reg[23][30]  ( .D(n368), .CK(clk), .RN(n2049), .Q(
        \register[23][30] ) );
  DFFRX1 \register_reg[23][29]  ( .D(n367), .CK(clk), .RN(n2048), .Q(
        \register[23][29] ) );
  DFFRX1 \register_reg[23][28]  ( .D(n366), .CK(clk), .RN(n2048), .Q(
        \register[23][28] ) );
  DFFRX1 \register_reg[23][27]  ( .D(n365), .CK(clk), .RN(n2048), .Q(
        \register[23][27] ) );
  DFFRX1 \register_reg[23][26]  ( .D(n364), .CK(clk), .RN(n2048), .Q(
        \register[23][26] ) );
  DFFRX1 \register_reg[23][25]  ( .D(n363), .CK(clk), .RN(n2048), .Q(
        \register[23][25] ) );
  DFFRX1 \register_reg[23][24]  ( .D(n362), .CK(clk), .RN(n2048), .Q(
        \register[23][24] ) );
  DFFRX1 \register_reg[23][23]  ( .D(n361), .CK(clk), .RN(n2048), .Q(
        \register[23][23] ) );
  DFFRX1 \register_reg[23][22]  ( .D(n360), .CK(clk), .RN(n2048), .Q(
        \register[23][22] ) );
  DFFRX1 \register_reg[23][21]  ( .D(n359), .CK(clk), .RN(n2048), .Q(
        \register[23][21] ) );
  DFFRX1 \register_reg[23][20]  ( .D(n358), .CK(clk), .RN(n2048), .Q(
        \register[23][20] ) );
  DFFRX1 \register_reg[23][19]  ( .D(n357), .CK(clk), .RN(n2048), .Q(
        \register[23][19] ) );
  DFFRX1 \register_reg[23][18]  ( .D(n356), .CK(clk), .RN(n2048), .Q(
        \register[23][18] ) );
  DFFRX1 \register_reg[23][17]  ( .D(n355), .CK(clk), .RN(n2048), .Q(
        \register[23][17] ) );
  DFFRX1 \register_reg[23][16]  ( .D(n354), .CK(clk), .RN(n2047), .Q(
        \register[23][16] ) );
  DFFRX1 \register_reg[23][15]  ( .D(n353), .CK(clk), .RN(n2047), .Q(
        \register[23][15] ) );
  DFFRX1 \register_reg[23][14]  ( .D(n352), .CK(clk), .RN(n2047), .Q(
        \register[23][14] ) );
  DFFRX1 \register_reg[23][13]  ( .D(n351), .CK(clk), .RN(n2047), .Q(
        \register[23][13] ) );
  DFFRX1 \register_reg[23][12]  ( .D(n350), .CK(clk), .RN(n2047), .Q(
        \register[23][12] ) );
  DFFRX1 \register_reg[23][11]  ( .D(n349), .CK(clk), .RN(n2047), .Q(
        \register[23][11] ) );
  DFFRX1 \register_reg[23][10]  ( .D(n348), .CK(clk), .RN(n2047), .Q(
        \register[23][10] ) );
  DFFRX1 \register_reg[23][9]  ( .D(n347), .CK(clk), .RN(n2047), .Q(
        \register[23][9] ) );
  DFFRX1 \register_reg[27][31]  ( .D(n241), .CK(clk), .RN(n2039), .Q(
        \register[27][31] ) );
  DFFRX1 \register_reg[27][30]  ( .D(n240), .CK(clk), .RN(n2039), .Q(
        \register[27][30] ) );
  DFFRX1 \register_reg[27][29]  ( .D(n239), .CK(clk), .RN(n2039), .Q(
        \register[27][29] ) );
  DFFRX1 \register_reg[27][28]  ( .D(n238), .CK(clk), .RN(n2039), .Q(
        \register[27][28] ) );
  DFFRX1 \register_reg[27][27]  ( .D(n237), .CK(clk), .RN(n2038), .Q(
        \register[27][27] ) );
  DFFRX1 \register_reg[27][26]  ( .D(n236), .CK(clk), .RN(n2038), .Q(
        \register[27][26] ) );
  DFFRX1 \register_reg[27][25]  ( .D(n235), .CK(clk), .RN(n2038), .Q(
        \register[27][25] ) );
  DFFRX1 \register_reg[27][24]  ( .D(n234), .CK(clk), .RN(n2038), .Q(
        \register[27][24] ) );
  DFFRX1 \register_reg[27][23]  ( .D(n233), .CK(clk), .RN(n2038), .Q(
        \register[27][23] ) );
  DFFRX1 \register_reg[27][22]  ( .D(n232), .CK(clk), .RN(n2038), .Q(
        \register[27][22] ) );
  DFFRX1 \register_reg[27][21]  ( .D(n231), .CK(clk), .RN(n2038), .Q(
        \register[27][21] ) );
  DFFRX1 \register_reg[27][20]  ( .D(n230), .CK(clk), .RN(n2038), .Q(
        \register[27][20] ) );
  DFFRX1 \register_reg[27][19]  ( .D(n229), .CK(clk), .RN(n2038), .Q(
        \register[27][19] ) );
  DFFRX1 \register_reg[27][18]  ( .D(n228), .CK(clk), .RN(n2038), .Q(
        \register[27][18] ) );
  DFFRX1 \register_reg[27][17]  ( .D(n227), .CK(clk), .RN(n2038), .Q(
        \register[27][17] ) );
  DFFRX1 \register_reg[27][16]  ( .D(n226), .CK(clk), .RN(n2038), .Q(
        \register[27][16] ) );
  DFFRX1 \register_reg[27][15]  ( .D(n225), .CK(clk), .RN(n2038), .Q(
        \register[27][15] ) );
  DFFRX1 \register_reg[27][14]  ( .D(n224), .CK(clk), .RN(n2037), .Q(
        \register[27][14] ) );
  DFFRX1 \register_reg[27][13]  ( .D(n223), .CK(clk), .RN(n2037), .Q(
        \register[27][13] ) );
  DFFRX1 \register_reg[27][12]  ( .D(n222), .CK(clk), .RN(n2037), .Q(
        \register[27][12] ) );
  DFFRX1 \register_reg[27][11]  ( .D(n221), .CK(clk), .RN(n2037), .Q(
        \register[27][11] ) );
  DFFRX1 \register_reg[27][10]  ( .D(n220), .CK(clk), .RN(n2037), .Q(
        \register[27][10] ) );
  DFFRX1 \register_reg[27][9]  ( .D(n219), .CK(clk), .RN(n2037), .Q(
        \register[27][9] ) );
  DFFRX1 \register_reg[31][31]  ( .D(n113), .CK(clk), .RN(n2029), .Q(
        \register[31][31] ) );
  DFFRX1 \register_reg[31][30]  ( .D(n112), .CK(clk), .RN(n2029), .Q(
        \register[31][30] ) );
  DFFRX1 \register_reg[31][29]  ( .D(n111), .CK(clk), .RN(n2029), .Q(
        \register[31][29] ) );
  DFFRX1 \register_reg[31][28]  ( .D(n110), .CK(clk), .RN(n2029), .Q(
        \register[31][28] ) );
  DFFRX1 \register_reg[31][27]  ( .D(n109), .CK(clk), .RN(n2029), .Q(
        \register[31][27] ) );
  DFFRX1 \register_reg[31][26]  ( .D(n108), .CK(clk), .RN(n2029), .Q(
        \register[31][26] ) );
  DFFRX1 \register_reg[31][25]  ( .D(n107), .CK(clk), .RN(n2028), .Q(
        \register[31][25] ) );
  DFFRX1 \register_reg[31][24]  ( .D(n106), .CK(clk), .RN(n2028), .Q(
        \register[31][24] ) );
  DFFRX1 \register_reg[31][23]  ( .D(n105), .CK(clk), .RN(n2028), .Q(
        \register[31][23] ) );
  DFFRX1 \register_reg[31][22]  ( .D(n104), .CK(clk), .RN(n2028), .Q(
        \register[31][22] ) );
  DFFRX1 \register_reg[31][21]  ( .D(n103), .CK(clk), .RN(n2028), .Q(
        \register[31][21] ) );
  DFFRX1 \register_reg[31][20]  ( .D(n102), .CK(clk), .RN(n2028), .Q(
        \register[31][20] ) );
  DFFRX1 \register_reg[31][19]  ( .D(n101), .CK(clk), .RN(n2028), .Q(
        \register[31][19] ) );
  DFFRX1 \register_reg[31][18]  ( .D(n100), .CK(clk), .RN(n2028), .Q(
        \register[31][18] ) );
  DFFRX1 \register_reg[31][17]  ( .D(n99), .CK(clk), .RN(n2028), .Q(
        \register[31][17] ) );
  DFFRX1 \register_reg[31][16]  ( .D(n98), .CK(clk), .RN(n2028), .Q(
        \register[31][16] ) );
  DFFRX1 \register_reg[31][15]  ( .D(n97), .CK(clk), .RN(n2028), .Q(
        \register[31][15] ) );
  DFFRX1 \register_reg[31][14]  ( .D(n96), .CK(clk), .RN(n2028), .Q(
        \register[31][14] ) );
  DFFRX1 \register_reg[31][13]  ( .D(n95), .CK(clk), .RN(n2028), .Q(
        \register[31][13] ) );
  DFFRX1 \register_reg[31][12]  ( .D(n94), .CK(clk), .RN(n2027), .Q(
        \register[31][12] ) );
  DFFRX1 \register_reg[31][11]  ( .D(n93), .CK(clk), .RN(n2027), .Q(
        \register[31][11] ) );
  DFFRX1 \register_reg[31][10]  ( .D(n92), .CK(clk), .RN(n2027), .Q(
        \register[31][10] ) );
  DFFRX1 \register_reg[31][9]  ( .D(n91), .CK(clk), .RN(n2027), .Q(
        \register[31][9] ) );
  DFFRX1 \register_reg[1][31]  ( .D(n1073), .CK(clk), .RN(n2103), .Q(
        \register[1][31] ) );
  DFFRX1 \register_reg[1][30]  ( .D(n1072), .CK(clk), .RN(n2103), .Q(
        \register[1][30] ) );
  DFFRX1 \register_reg[1][29]  ( .D(n1071), .CK(clk), .RN(n2103), .Q(
        \register[1][29] ) );
  DFFRX1 \register_reg[1][28]  ( .D(n1070), .CK(clk), .RN(n2103), .Q(
        \register[1][28] ) );
  DFFRX1 \register_reg[1][27]  ( .D(n1069), .CK(clk), .RN(n2102), .Q(
        \register[1][27] ) );
  DFFRX1 \register_reg[1][26]  ( .D(n1068), .CK(clk), .RN(n2102), .Q(
        \register[1][26] ) );
  DFFRX1 \register_reg[1][25]  ( .D(n1067), .CK(clk), .RN(n2102), .Q(
        \register[1][25] ) );
  DFFRX1 \register_reg[1][24]  ( .D(n1066), .CK(clk), .RN(n2102), .Q(
        \register[1][24] ) );
  DFFRX1 \register_reg[1][23]  ( .D(n1065), .CK(clk), .RN(n2102), .Q(
        \register[1][23] ) );
  DFFRX1 \register_reg[1][22]  ( .D(n1064), .CK(clk), .RN(n2102), .Q(
        \register[1][22] ) );
  DFFRX1 \register_reg[1][21]  ( .D(n1063), .CK(clk), .RN(n2102), .Q(
        \register[1][21] ) );
  DFFRX1 \register_reg[1][20]  ( .D(n1062), .CK(clk), .RN(n2102), .Q(
        \register[1][20] ) );
  DFFRX1 \register_reg[1][19]  ( .D(n1061), .CK(clk), .RN(n2102), .Q(
        \register[1][19] ) );
  DFFRX1 \register_reg[1][18]  ( .D(n1060), .CK(clk), .RN(n2102), .Q(
        \register[1][18] ) );
  DFFRX1 \register_reg[1][17]  ( .D(n1059), .CK(clk), .RN(n2102), .Q(
        \register[1][17] ) );
  DFFRX1 \register_reg[1][16]  ( .D(n1058), .CK(clk), .RN(n2102), .Q(
        \register[1][16] ) );
  DFFRX1 \register_reg[1][15]  ( .D(n1057), .CK(clk), .RN(n2102), .Q(
        \register[1][15] ) );
  DFFRX1 \register_reg[1][14]  ( .D(n1056), .CK(clk), .RN(n2101), .Q(
        \register[1][14] ) );
  DFFRX1 \register_reg[1][13]  ( .D(n1055), .CK(clk), .RN(n2101), .Q(
        \register[1][13] ) );
  DFFRX1 \register_reg[1][12]  ( .D(n1054), .CK(clk), .RN(n2101), .Q(
        \register[1][12] ) );
  DFFRX1 \register_reg[1][11]  ( .D(n1053), .CK(clk), .RN(n2101), .Q(
        \register[1][11] ) );
  DFFRX1 \register_reg[1][10]  ( .D(n1052), .CK(clk), .RN(n2101), .Q(
        \register[1][10] ) );
  DFFRX1 \register_reg[1][9]  ( .D(n1051), .CK(clk), .RN(n2101), .Q(
        \register[1][9] ) );
  DFFRX1 \register_reg[5][31]  ( .D(n945), .CK(clk), .RN(n2093), .Q(
        \register[5][31] ) );
  DFFRX1 \register_reg[5][30]  ( .D(n944), .CK(clk), .RN(n2093), .Q(
        \register[5][30] ) );
  DFFRX1 \register_reg[5][29]  ( .D(n943), .CK(clk), .RN(n2093), .Q(
        \register[5][29] ) );
  DFFRX1 \register_reg[5][28]  ( .D(n942), .CK(clk), .RN(n2093), .Q(
        \register[5][28] ) );
  DFFRX1 \register_reg[5][27]  ( .D(n941), .CK(clk), .RN(n2093), .Q(
        \register[5][27] ) );
  DFFRX1 \register_reg[5][26]  ( .D(n940), .CK(clk), .RN(n2093), .Q(
        \register[5][26] ) );
  DFFRX1 \register_reg[5][25]  ( .D(n939), .CK(clk), .RN(n2092), .Q(
        \register[5][25] ) );
  DFFRX1 \register_reg[5][24]  ( .D(n938), .CK(clk), .RN(n2092), .Q(
        \register[5][24] ) );
  DFFRX1 \register_reg[5][23]  ( .D(n937), .CK(clk), .RN(n2092), .Q(
        \register[5][23] ) );
  DFFRX1 \register_reg[5][22]  ( .D(n936), .CK(clk), .RN(n2092), .Q(
        \register[5][22] ) );
  DFFRX1 \register_reg[5][21]  ( .D(n935), .CK(clk), .RN(n2092), .Q(
        \register[5][21] ) );
  DFFRX1 \register_reg[5][20]  ( .D(n934), .CK(clk), .RN(n2092), .Q(
        \register[5][20] ) );
  DFFRX1 \register_reg[5][19]  ( .D(n933), .CK(clk), .RN(n2092), .Q(
        \register[5][19] ) );
  DFFRX1 \register_reg[5][18]  ( .D(n932), .CK(clk), .RN(n2092), .Q(
        \register[5][18] ) );
  DFFRX1 \register_reg[5][17]  ( .D(n931), .CK(clk), .RN(n2092), .Q(
        \register[5][17] ) );
  DFFRX1 \register_reg[5][16]  ( .D(n930), .CK(clk), .RN(n2092), .Q(
        \register[5][16] ) );
  DFFRX1 \register_reg[5][15]  ( .D(n929), .CK(clk), .RN(n2092), .Q(
        \register[5][15] ) );
  DFFRX1 \register_reg[5][14]  ( .D(n928), .CK(clk), .RN(n2092), .Q(
        \register[5][14] ) );
  DFFRX1 \register_reg[5][13]  ( .D(n927), .CK(clk), .RN(n2092), .Q(
        \register[5][13] ) );
  DFFRX1 \register_reg[5][12]  ( .D(n926), .CK(clk), .RN(n2091), .Q(
        \register[5][12] ) );
  DFFRX1 \register_reg[5][11]  ( .D(n925), .CK(clk), .RN(n2091), .Q(
        \register[5][11] ) );
  DFFRX1 \register_reg[5][10]  ( .D(n924), .CK(clk), .RN(n2091), .Q(
        \register[5][10] ) );
  DFFRX1 \register_reg[5][9]  ( .D(n923), .CK(clk), .RN(n2091), .Q(
        \register[5][9] ) );
  DFFRX1 \register_reg[9][31]  ( .D(n817), .CK(clk), .RN(n2083), .Q(
        \register[9][31] ) );
  DFFRX1 \register_reg[9][30]  ( .D(n816), .CK(clk), .RN(n2083), .Q(
        \register[9][30] ) );
  DFFRX1 \register_reg[9][29]  ( .D(n815), .CK(clk), .RN(n2083), .Q(
        \register[9][29] ) );
  DFFRX1 \register_reg[9][28]  ( .D(n814), .CK(clk), .RN(n2083), .Q(
        \register[9][28] ) );
  DFFRX1 \register_reg[9][27]  ( .D(n813), .CK(clk), .RN(n2083), .Q(
        \register[9][27] ) );
  DFFRX1 \register_reg[9][26]  ( .D(n812), .CK(clk), .RN(n2083), .Q(
        \register[9][26] ) );
  DFFRX1 \register_reg[9][25]  ( .D(n811), .CK(clk), .RN(n2083), .Q(
        \register[9][25] ) );
  DFFRX1 \register_reg[9][24]  ( .D(n810), .CK(clk), .RN(n2083), .Q(
        \register[9][24] ) );
  DFFRX1 \register_reg[9][23]  ( .D(n809), .CK(clk), .RN(n2082), .Q(
        \register[9][23] ) );
  DFFRX1 \register_reg[9][22]  ( .D(n808), .CK(clk), .RN(n2082), .Q(
        \register[9][22] ) );
  DFFRX1 \register_reg[9][21]  ( .D(n807), .CK(clk), .RN(n2082), .Q(
        \register[9][21] ) );
  DFFRX1 \register_reg[9][20]  ( .D(n806), .CK(clk), .RN(n2082), .Q(
        \register[9][20] ) );
  DFFRX1 \register_reg[9][19]  ( .D(n805), .CK(clk), .RN(n2082), .Q(
        \register[9][19] ) );
  DFFRX1 \register_reg[9][18]  ( .D(n804), .CK(clk), .RN(n2082), .Q(
        \register[9][18] ) );
  DFFRX1 \register_reg[9][17]  ( .D(n803), .CK(clk), .RN(n2082), .Q(
        \register[9][17] ) );
  DFFRX1 \register_reg[9][16]  ( .D(n802), .CK(clk), .RN(n2082), .Q(
        \register[9][16] ) );
  DFFRX1 \register_reg[9][15]  ( .D(n801), .CK(clk), .RN(n2082), .Q(
        \register[9][15] ) );
  DFFRX1 \register_reg[9][14]  ( .D(n800), .CK(clk), .RN(n2082), .Q(
        \register[9][14] ) );
  DFFRX1 \register_reg[9][13]  ( .D(n799), .CK(clk), .RN(n2082), .Q(
        \register[9][13] ) );
  DFFRX1 \register_reg[9][12]  ( .D(n798), .CK(clk), .RN(n2082), .Q(
        \register[9][12] ) );
  DFFRX1 \register_reg[9][11]  ( .D(n797), .CK(clk), .RN(n2082), .Q(
        \register[9][11] ) );
  DFFRX1 \register_reg[9][10]  ( .D(n796), .CK(clk), .RN(n2081), .Q(
        \register[9][10] ) );
  DFFRX1 \register_reg[9][9]  ( .D(n795), .CK(clk), .RN(n2081), .Q(
        \register[9][9] ) );
  DFFRX1 \register_reg[13][31]  ( .D(n689), .CK(clk), .RN(n2073), .Q(
        \register[13][31] ) );
  DFFRX1 \register_reg[13][30]  ( .D(n688), .CK(clk), .RN(n2073), .Q(
        \register[13][30] ) );
  DFFRX1 \register_reg[13][29]  ( .D(n687), .CK(clk), .RN(n2073), .Q(
        \register[13][29] ) );
  DFFRX1 \register_reg[13][28]  ( .D(n686), .CK(clk), .RN(n2073), .Q(
        \register[13][28] ) );
  DFFRX1 \register_reg[13][27]  ( .D(n685), .CK(clk), .RN(n2073), .Q(
        \register[13][27] ) );
  DFFRX1 \register_reg[13][26]  ( .D(n684), .CK(clk), .RN(n2073), .Q(
        \register[13][26] ) );
  DFFRX1 \register_reg[13][25]  ( .D(n683), .CK(clk), .RN(n2073), .Q(
        \register[13][25] ) );
  DFFRX1 \register_reg[13][24]  ( .D(n682), .CK(clk), .RN(n2073), .Q(
        \register[13][24] ) );
  DFFRX1 \register_reg[13][23]  ( .D(n681), .CK(clk), .RN(n2073), .Q(
        \register[13][23] ) );
  DFFRX1 \register_reg[13][22]  ( .D(n680), .CK(clk), .RN(n2073), .Q(
        \register[13][22] ) );
  DFFRX1 \register_reg[13][21]  ( .D(n679), .CK(clk), .RN(n2072), .Q(
        \register[13][21] ) );
  DFFRX1 \register_reg[13][20]  ( .D(n678), .CK(clk), .RN(n2072), .Q(
        \register[13][20] ) );
  DFFRX1 \register_reg[13][19]  ( .D(n677), .CK(clk), .RN(n2072), .Q(
        \register[13][19] ) );
  DFFRX1 \register_reg[13][18]  ( .D(n676), .CK(clk), .RN(n2072), .Q(
        \register[13][18] ) );
  DFFRX1 \register_reg[13][17]  ( .D(n675), .CK(clk), .RN(n2072), .Q(
        \register[13][17] ) );
  DFFRX1 \register_reg[13][16]  ( .D(n674), .CK(clk), .RN(n2072), .Q(
        \register[13][16] ) );
  DFFRX1 \register_reg[13][15]  ( .D(n673), .CK(clk), .RN(n2072), .Q(
        \register[13][15] ) );
  DFFRX1 \register_reg[13][14]  ( .D(n672), .CK(clk), .RN(n2072), .Q(
        \register[13][14] ) );
  DFFRX1 \register_reg[13][13]  ( .D(n671), .CK(clk), .RN(n2072), .Q(
        \register[13][13] ) );
  DFFRX1 \register_reg[13][12]  ( .D(n670), .CK(clk), .RN(n2072), .Q(
        \register[13][12] ) );
  DFFRX1 \register_reg[13][11]  ( .D(n669), .CK(clk), .RN(n2072), .Q(
        \register[13][11] ) );
  DFFRX1 \register_reg[13][10]  ( .D(n668), .CK(clk), .RN(n2072), .Q(
        \register[13][10] ) );
  DFFRX1 \register_reg[13][9]  ( .D(n667), .CK(clk), .RN(n2072), .Q(
        \register[13][9] ) );
  DFFRX1 \register_reg[17][31]  ( .D(n561), .CK(clk), .RN(n2063), .Q(
        \register[17][31] ) );
  DFFRX1 \register_reg[17][30]  ( .D(n560), .CK(clk), .RN(n2063), .Q(
        \register[17][30] ) );
  DFFRX1 \register_reg[17][29]  ( .D(n559), .CK(clk), .RN(n2063), .Q(
        \register[17][29] ) );
  DFFRX1 \register_reg[17][28]  ( .D(n558), .CK(clk), .RN(n2063), .Q(
        \register[17][28] ) );
  DFFRX1 \register_reg[17][27]  ( .D(n557), .CK(clk), .RN(n2063), .Q(
        \register[17][27] ) );
  DFFRX1 \register_reg[17][26]  ( .D(n556), .CK(clk), .RN(n2063), .Q(
        \register[17][26] ) );
  DFFRX1 \register_reg[17][25]  ( .D(n555), .CK(clk), .RN(n2063), .Q(
        \register[17][25] ) );
  DFFRX1 \register_reg[17][24]  ( .D(n554), .CK(clk), .RN(n2063), .Q(
        \register[17][24] ) );
  DFFRX1 \register_reg[17][23]  ( .D(n553), .CK(clk), .RN(n2063), .Q(
        \register[17][23] ) );
  DFFRX1 \register_reg[17][22]  ( .D(n552), .CK(clk), .RN(n2063), .Q(
        \register[17][22] ) );
  DFFRX1 \register_reg[17][21]  ( .D(n551), .CK(clk), .RN(n2063), .Q(
        \register[17][21] ) );
  DFFRX1 \register_reg[17][20]  ( .D(n550), .CK(clk), .RN(n2063), .Q(
        \register[17][20] ) );
  DFFRX1 \register_reg[17][19]  ( .D(n549), .CK(clk), .RN(n2062), .Q(
        \register[17][19] ) );
  DFFRX1 \register_reg[17][18]  ( .D(n548), .CK(clk), .RN(n2062), .Q(
        \register[17][18] ) );
  DFFRX1 \register_reg[17][17]  ( .D(n547), .CK(clk), .RN(n2062), .Q(
        \register[17][17] ) );
  DFFRX1 \register_reg[17][16]  ( .D(n546), .CK(clk), .RN(n2062), .Q(
        \register[17][16] ) );
  DFFRX1 \register_reg[17][15]  ( .D(n545), .CK(clk), .RN(n2062), .Q(
        \register[17][15] ) );
  DFFRX1 \register_reg[17][14]  ( .D(n544), .CK(clk), .RN(n2062), .Q(
        \register[17][14] ) );
  DFFRX1 \register_reg[17][13]  ( .D(n543), .CK(clk), .RN(n2062), .Q(
        \register[17][13] ) );
  DFFRX1 \register_reg[17][12]  ( .D(n542), .CK(clk), .RN(n2062), .Q(
        \register[17][12] ) );
  DFFRX1 \register_reg[17][11]  ( .D(n541), .CK(clk), .RN(n2062), .Q(
        \register[17][11] ) );
  DFFRX1 \register_reg[17][10]  ( .D(n540), .CK(clk), .RN(n2062), .Q(
        \register[17][10] ) );
  DFFRX1 \register_reg[17][9]  ( .D(n539), .CK(clk), .RN(n2062), .Q(
        \register[17][9] ) );
  DFFRX1 \register_reg[21][31]  ( .D(n433), .CK(clk), .RN(n2054), .Q(
        \register[21][31] ) );
  DFFRX1 \register_reg[21][30]  ( .D(n432), .CK(clk), .RN(n2053), .Q(
        \register[21][30] ) );
  DFFRX1 \register_reg[21][29]  ( .D(n431), .CK(clk), .RN(n2053), .Q(
        \register[21][29] ) );
  DFFRX1 \register_reg[21][28]  ( .D(n430), .CK(clk), .RN(n2053), .Q(
        \register[21][28] ) );
  DFFRX1 \register_reg[21][27]  ( .D(n429), .CK(clk), .RN(n2053), .Q(
        \register[21][27] ) );
  DFFRX1 \register_reg[21][26]  ( .D(n428), .CK(clk), .RN(n2053), .Q(
        \register[21][26] ) );
  DFFRX1 \register_reg[21][25]  ( .D(n427), .CK(clk), .RN(n2053), .Q(
        \register[21][25] ) );
  DFFRX1 \register_reg[21][24]  ( .D(n426), .CK(clk), .RN(n2053), .Q(
        \register[21][24] ) );
  DFFRX1 \register_reg[21][23]  ( .D(n425), .CK(clk), .RN(n2053), .Q(
        \register[21][23] ) );
  DFFRX1 \register_reg[21][22]  ( .D(n424), .CK(clk), .RN(n2053), .Q(
        \register[21][22] ) );
  DFFRX1 \register_reg[21][21]  ( .D(n423), .CK(clk), .RN(n2053), .Q(
        \register[21][21] ) );
  DFFRX1 \register_reg[21][20]  ( .D(n422), .CK(clk), .RN(n2053), .Q(
        \register[21][20] ) );
  DFFRX1 \register_reg[21][19]  ( .D(n421), .CK(clk), .RN(n2053), .Q(
        \register[21][19] ) );
  DFFRX1 \register_reg[21][18]  ( .D(n420), .CK(clk), .RN(n2053), .Q(
        \register[21][18] ) );
  DFFRX1 \register_reg[21][17]  ( .D(n419), .CK(clk), .RN(n2052), .Q(
        \register[21][17] ) );
  DFFRX1 \register_reg[21][16]  ( .D(n418), .CK(clk), .RN(n2052), .Q(
        \register[21][16] ) );
  DFFRX1 \register_reg[21][15]  ( .D(n417), .CK(clk), .RN(n2052), .Q(
        \register[21][15] ) );
  DFFRX1 \register_reg[21][14]  ( .D(n416), .CK(clk), .RN(n2052), .Q(
        \register[21][14] ) );
  DFFRX1 \register_reg[21][13]  ( .D(n415), .CK(clk), .RN(n2052), .Q(
        \register[21][13] ) );
  DFFRX1 \register_reg[21][12]  ( .D(n414), .CK(clk), .RN(n2052), .Q(
        \register[21][12] ) );
  DFFRX1 \register_reg[21][11]  ( .D(n413), .CK(clk), .RN(n2052), .Q(
        \register[21][11] ) );
  DFFRX1 \register_reg[21][10]  ( .D(n412), .CK(clk), .RN(n2052), .Q(
        \register[21][10] ) );
  DFFRX1 \register_reg[21][9]  ( .D(n411), .CK(clk), .RN(n2052), .Q(
        \register[21][9] ) );
  DFFRX1 \register_reg[25][31]  ( .D(n305), .CK(clk), .RN(n2044), .Q(
        \register[25][31] ) );
  DFFRX1 \register_reg[25][30]  ( .D(n304), .CK(clk), .RN(n2044), .Q(
        \register[25][30] ) );
  DFFRX1 \register_reg[25][29]  ( .D(n303), .CK(clk), .RN(n2044), .Q(
        \register[25][29] ) );
  DFFRX1 \register_reg[25][28]  ( .D(n302), .CK(clk), .RN(n2043), .Q(
        \register[25][28] ) );
  DFFRX1 \register_reg[25][27]  ( .D(n301), .CK(clk), .RN(n2043), .Q(
        \register[25][27] ) );
  DFFRX1 \register_reg[25][26]  ( .D(n300), .CK(clk), .RN(n2043), .Q(
        \register[25][26] ) );
  DFFRX1 \register_reg[25][25]  ( .D(n299), .CK(clk), .RN(n2043), .Q(
        \register[25][25] ) );
  DFFRX1 \register_reg[25][24]  ( .D(n298), .CK(clk), .RN(n2043), .Q(
        \register[25][24] ) );
  DFFRX1 \register_reg[25][23]  ( .D(n297), .CK(clk), .RN(n2043), .Q(
        \register[25][23] ) );
  DFFRX1 \register_reg[25][22]  ( .D(n296), .CK(clk), .RN(n2043), .Q(
        \register[25][22] ) );
  DFFRX1 \register_reg[25][21]  ( .D(n295), .CK(clk), .RN(n2043), .Q(
        \register[25][21] ) );
  DFFRX1 \register_reg[25][20]  ( .D(n294), .CK(clk), .RN(n2043), .Q(
        \register[25][20] ) );
  DFFRX1 \register_reg[25][19]  ( .D(n293), .CK(clk), .RN(n2043), .Q(
        \register[25][19] ) );
  DFFRX1 \register_reg[25][18]  ( .D(n292), .CK(clk), .RN(n2043), .Q(
        \register[25][18] ) );
  DFFRX1 \register_reg[25][17]  ( .D(n291), .CK(clk), .RN(n2043), .Q(
        \register[25][17] ) );
  DFFRX1 \register_reg[25][16]  ( .D(n290), .CK(clk), .RN(n2043), .Q(
        \register[25][16] ) );
  DFFRX1 \register_reg[25][15]  ( .D(n289), .CK(clk), .RN(n2042), .Q(
        \register[25][15] ) );
  DFFRX1 \register_reg[25][14]  ( .D(n288), .CK(clk), .RN(n2042), .Q(
        \register[25][14] ) );
  DFFRX1 \register_reg[25][13]  ( .D(n287), .CK(clk), .RN(n2042), .Q(
        \register[25][13] ) );
  DFFRX1 \register_reg[25][12]  ( .D(n286), .CK(clk), .RN(n2042), .Q(
        \register[25][12] ) );
  DFFRX1 \register_reg[25][11]  ( .D(n285), .CK(clk), .RN(n2042), .Q(
        \register[25][11] ) );
  DFFRX1 \register_reg[25][10]  ( .D(n284), .CK(clk), .RN(n2042), .Q(
        \register[25][10] ) );
  DFFRX1 \register_reg[25][9]  ( .D(n283), .CK(clk), .RN(n2042), .Q(
        \register[25][9] ) );
  DFFRX1 \register_reg[29][31]  ( .D(n177), .CK(clk), .RN(n2034), .Q(
        \register[29][31] ) );
  DFFRX1 \register_reg[29][30]  ( .D(n176), .CK(clk), .RN(n2034), .Q(
        \register[29][30] ) );
  DFFRX1 \register_reg[29][29]  ( .D(n175), .CK(clk), .RN(n2034), .Q(
        \register[29][29] ) );
  DFFRX1 \register_reg[29][28]  ( .D(n174), .CK(clk), .RN(n2034), .Q(
        \register[29][28] ) );
  DFFRX1 \register_reg[29][27]  ( .D(n173), .CK(clk), .RN(n2034), .Q(
        \register[29][27] ) );
  DFFRX1 \register_reg[29][26]  ( .D(n172), .CK(clk), .RN(n2033), .Q(
        \register[29][26] ) );
  DFFRX1 \register_reg[29][25]  ( .D(n171), .CK(clk), .RN(n2033), .Q(
        \register[29][25] ) );
  DFFRX1 \register_reg[29][24]  ( .D(n170), .CK(clk), .RN(n2033), .Q(
        \register[29][24] ) );
  DFFRX1 \register_reg[29][23]  ( .D(n169), .CK(clk), .RN(n2033), .Q(
        \register[29][23] ) );
  DFFRX1 \register_reg[29][22]  ( .D(n168), .CK(clk), .RN(n2033), .Q(
        \register[29][22] ) );
  DFFRX1 \register_reg[29][21]  ( .D(n167), .CK(clk), .RN(n2033), .Q(
        \register[29][21] ) );
  DFFRX1 \register_reg[29][20]  ( .D(n166), .CK(clk), .RN(n2033), .Q(
        \register[29][20] ) );
  DFFRX1 \register_reg[29][19]  ( .D(n165), .CK(clk), .RN(n2033), .Q(
        \register[29][19] ) );
  DFFRX1 \register_reg[29][18]  ( .D(n164), .CK(clk), .RN(n2033), .Q(
        \register[29][18] ) );
  DFFRX1 \register_reg[29][17]  ( .D(n163), .CK(clk), .RN(n2033), .Q(
        \register[29][17] ) );
  DFFRX1 \register_reg[29][16]  ( .D(n162), .CK(clk), .RN(n2033), .Q(
        \register[29][16] ) );
  DFFRX1 \register_reg[29][15]  ( .D(n161), .CK(clk), .RN(n2033), .Q(
        \register[29][15] ) );
  DFFRX1 \register_reg[29][14]  ( .D(n160), .CK(clk), .RN(n2033), .Q(
        \register[29][14] ) );
  DFFRX1 \register_reg[29][13]  ( .D(n159), .CK(clk), .RN(n2032), .Q(
        \register[29][13] ) );
  DFFRX1 \register_reg[29][12]  ( .D(n158), .CK(clk), .RN(n2032), .Q(
        \register[29][12] ) );
  DFFRX1 \register_reg[29][11]  ( .D(n157), .CK(clk), .RN(n2032), .Q(
        \register[29][11] ) );
  DFFRX1 \register_reg[29][10]  ( .D(n156), .CK(clk), .RN(n2032), .Q(
        \register[29][10] ) );
  DFFRX1 \register_reg[29][9]  ( .D(n155), .CK(clk), .RN(n2032), .Q(
        \register[29][9] ) );
  DFFRX1 \register_reg[0][31]  ( .D(n1105), .CK(clk), .RN(n2105), .Q(
        \register[0][31] ) );
  DFFRX1 \register_reg[0][30]  ( .D(n1104), .CK(clk), .RN(n2105), .Q(
        \register[0][30] ) );
  DFFRX1 \register_reg[0][29]  ( .D(n1103), .CK(clk), .RN(n2105), .Q(
        \register[0][29] ) );
  DFFRX1 \register_reg[0][28]  ( .D(n1102), .CK(clk), .RN(n2105), .Q(
        \register[0][28] ) );
  DFFRX1 \register_reg[0][27]  ( .D(n1101), .CK(clk), .RN(n2105), .Q(
        \register[0][27] ) );
  DFFRX1 \register_reg[0][26]  ( .D(n1100), .CK(clk), .RN(n2105), .Q(
        \register[0][26] ) );
  DFFRX1 \register_reg[0][25]  ( .D(n1099), .CK(clk), .RN(n2105), .Q(
        \register[0][25] ) );
  DFFRX1 \register_reg[0][24]  ( .D(n1098), .CK(clk), .RN(n2105), .Q(
        \register[0][24] ) );
  DFFRX1 \register_reg[0][23]  ( .D(n1097), .CK(clk), .RN(n2105), .Q(
        \register[0][23] ) );
  DFFRX1 \register_reg[0][22]  ( .D(n1096), .CK(clk), .RN(n2105), .Q(
        \register[0][22] ) );
  DFFRX1 \register_reg[0][21]  ( .D(n1095), .CK(clk), .RN(n2104), .Q(
        \register[0][21] ) );
  DFFRX1 \register_reg[0][20]  ( .D(n1094), .CK(clk), .RN(n2104), .Q(
        \register[0][20] ) );
  DFFRX1 \register_reg[0][19]  ( .D(n1093), .CK(clk), .RN(n2104), .Q(
        \register[0][19] ) );
  DFFRX1 \register_reg[0][18]  ( .D(n1092), .CK(clk), .RN(n2104), .Q(
        \register[0][18] ) );
  DFFRX1 \register_reg[0][17]  ( .D(n1091), .CK(clk), .RN(n2104), .Q(
        \register[0][17] ) );
  DFFRX1 \register_reg[0][16]  ( .D(n1090), .CK(clk), .RN(n2104), .Q(
        \register[0][16] ) );
  DFFRX1 \register_reg[0][15]  ( .D(n1089), .CK(clk), .RN(n2104), .Q(
        \register[0][15] ) );
  DFFRX1 \register_reg[0][14]  ( .D(n1088), .CK(clk), .RN(n2104), .Q(
        \register[0][14] ) );
  DFFRX1 \register_reg[0][13]  ( .D(n1087), .CK(clk), .RN(n2104), .Q(
        \register[0][13] ) );
  DFFRX1 \register_reg[0][12]  ( .D(n1086), .CK(clk), .RN(n2104), .Q(
        \register[0][12] ) );
  DFFRX1 \register_reg[0][11]  ( .D(n1085), .CK(clk), .RN(n2104), .Q(
        \register[0][11] ) );
  DFFRX1 \register_reg[0][10]  ( .D(n1084), .CK(clk), .RN(n2104), .Q(
        \register[0][10] ) );
  DFFRX1 \register_reg[0][9]  ( .D(n1083), .CK(clk), .RN(n2104), .Q(
        \register[0][9] ) );
  DFFRX1 \register_reg[4][31]  ( .D(n977), .CK(clk), .RN(n2095), .Q(
        \register[4][31] ) );
  DFFRX1 \register_reg[4][30]  ( .D(n976), .CK(clk), .RN(n2095), .Q(
        \register[4][30] ) );
  DFFRX1 \register_reg[4][29]  ( .D(n975), .CK(clk), .RN(n2095), .Q(
        \register[4][29] ) );
  DFFRX1 \register_reg[4][28]  ( .D(n974), .CK(clk), .RN(n2095), .Q(
        \register[4][28] ) );
  DFFRX1 \register_reg[4][27]  ( .D(n973), .CK(clk), .RN(n2095), .Q(
        \register[4][27] ) );
  DFFRX1 \register_reg[4][26]  ( .D(n972), .CK(clk), .RN(n2095), .Q(
        \register[4][26] ) );
  DFFRX1 \register_reg[4][25]  ( .D(n971), .CK(clk), .RN(n2095), .Q(
        \register[4][25] ) );
  DFFRX1 \register_reg[4][24]  ( .D(n970), .CK(clk), .RN(n2095), .Q(
        \register[4][24] ) );
  DFFRX1 \register_reg[4][23]  ( .D(n969), .CK(clk), .RN(n2095), .Q(
        \register[4][23] ) );
  DFFRX1 \register_reg[4][22]  ( .D(n968), .CK(clk), .RN(n2095), .Q(
        \register[4][22] ) );
  DFFRX1 \register_reg[4][21]  ( .D(n967), .CK(clk), .RN(n2095), .Q(
        \register[4][21] ) );
  DFFRX1 \register_reg[4][20]  ( .D(n966), .CK(clk), .RN(n2095), .Q(
        \register[4][20] ) );
  DFFRX1 \register_reg[4][19]  ( .D(n965), .CK(clk), .RN(n2094), .Q(
        \register[4][19] ) );
  DFFRX1 \register_reg[4][18]  ( .D(n964), .CK(clk), .RN(n2094), .Q(
        \register[4][18] ) );
  DFFRX1 \register_reg[4][17]  ( .D(n963), .CK(clk), .RN(n2094), .Q(
        \register[4][17] ) );
  DFFRX1 \register_reg[4][16]  ( .D(n962), .CK(clk), .RN(n2094), .Q(
        \register[4][16] ) );
  DFFRX1 \register_reg[4][15]  ( .D(n961), .CK(clk), .RN(n2094), .Q(
        \register[4][15] ) );
  DFFRX1 \register_reg[4][14]  ( .D(n960), .CK(clk), .RN(n2094), .Q(
        \register[4][14] ) );
  DFFRX1 \register_reg[4][13]  ( .D(n959), .CK(clk), .RN(n2094), .Q(
        \register[4][13] ) );
  DFFRX1 \register_reg[4][12]  ( .D(n958), .CK(clk), .RN(n2094), .Q(
        \register[4][12] ) );
  DFFRX1 \register_reg[4][11]  ( .D(n957), .CK(clk), .RN(n2094), .Q(
        \register[4][11] ) );
  DFFRX1 \register_reg[4][10]  ( .D(n956), .CK(clk), .RN(n2094), .Q(
        \register[4][10] ) );
  DFFRX1 \register_reg[4][9]  ( .D(n955), .CK(clk), .RN(n2094), .Q(
        \register[4][9] ) );
  DFFRX1 \register_reg[8][31]  ( .D(n849), .CK(clk), .RN(n2086), .Q(
        \register[8][31] ) );
  DFFRX1 \register_reg[8][30]  ( .D(n848), .CK(clk), .RN(n2085), .Q(
        \register[8][30] ) );
  DFFRX1 \register_reg[8][29]  ( .D(n847), .CK(clk), .RN(n2085), .Q(
        \register[8][29] ) );
  DFFRX1 \register_reg[8][28]  ( .D(n846), .CK(clk), .RN(n2085), .Q(
        \register[8][28] ) );
  DFFRX1 \register_reg[8][27]  ( .D(n845), .CK(clk), .RN(n2085), .Q(
        \register[8][27] ) );
  DFFRX1 \register_reg[8][26]  ( .D(n844), .CK(clk), .RN(n2085), .Q(
        \register[8][26] ) );
  DFFRX1 \register_reg[8][25]  ( .D(n843), .CK(clk), .RN(n2085), .Q(
        \register[8][25] ) );
  DFFRX1 \register_reg[8][24]  ( .D(n842), .CK(clk), .RN(n2085), .Q(
        \register[8][24] ) );
  DFFRX1 \register_reg[8][23]  ( .D(n841), .CK(clk), .RN(n2085), .Q(
        \register[8][23] ) );
  DFFRX1 \register_reg[8][22]  ( .D(n840), .CK(clk), .RN(n2085), .Q(
        \register[8][22] ) );
  DFFRX1 \register_reg[8][21]  ( .D(n839), .CK(clk), .RN(n2085), .Q(
        \register[8][21] ) );
  DFFRX1 \register_reg[8][20]  ( .D(n838), .CK(clk), .RN(n2085), .Q(
        \register[8][20] ) );
  DFFRX1 \register_reg[8][19]  ( .D(n837), .CK(clk), .RN(n2085), .Q(
        \register[8][19] ) );
  DFFRX1 \register_reg[8][18]  ( .D(n836), .CK(clk), .RN(n2085), .Q(
        \register[8][18] ) );
  DFFRX1 \register_reg[8][17]  ( .D(n835), .CK(clk), .RN(n2084), .Q(
        \register[8][17] ) );
  DFFRX1 \register_reg[8][16]  ( .D(n834), .CK(clk), .RN(n2084), .Q(
        \register[8][16] ) );
  DFFRX1 \register_reg[8][15]  ( .D(n833), .CK(clk), .RN(n2084), .Q(
        \register[8][15] ) );
  DFFRX1 \register_reg[8][14]  ( .D(n832), .CK(clk), .RN(n2084), .Q(
        \register[8][14] ) );
  DFFRX1 \register_reg[8][13]  ( .D(n831), .CK(clk), .RN(n2084), .Q(
        \register[8][13] ) );
  DFFRX1 \register_reg[8][12]  ( .D(n830), .CK(clk), .RN(n2084), .Q(
        \register[8][12] ) );
  DFFRX1 \register_reg[8][11]  ( .D(n829), .CK(clk), .RN(n2084), .Q(
        \register[8][11] ) );
  DFFRX1 \register_reg[8][10]  ( .D(n828), .CK(clk), .RN(n2084), .Q(
        \register[8][10] ) );
  DFFRX1 \register_reg[8][9]  ( .D(n827), .CK(clk), .RN(n2084), .Q(
        \register[8][9] ) );
  DFFRX1 \register_reg[12][31]  ( .D(n721), .CK(clk), .RN(n2076), .Q(
        \register[12][31] ) );
  DFFRX1 \register_reg[12][30]  ( .D(n720), .CK(clk), .RN(n2076), .Q(
        \register[12][30] ) );
  DFFRX1 \register_reg[12][29]  ( .D(n719), .CK(clk), .RN(n2076), .Q(
        \register[12][29] ) );
  DFFRX1 \register_reg[12][28]  ( .D(n718), .CK(clk), .RN(n2075), .Q(
        \register[12][28] ) );
  DFFRX1 \register_reg[12][27]  ( .D(n717), .CK(clk), .RN(n2075), .Q(
        \register[12][27] ) );
  DFFRX1 \register_reg[12][26]  ( .D(n716), .CK(clk), .RN(n2075), .Q(
        \register[12][26] ) );
  DFFRX1 \register_reg[12][25]  ( .D(n715), .CK(clk), .RN(n2075), .Q(
        \register[12][25] ) );
  DFFRX1 \register_reg[12][24]  ( .D(n714), .CK(clk), .RN(n2075), .Q(
        \register[12][24] ) );
  DFFRX1 \register_reg[12][23]  ( .D(n713), .CK(clk), .RN(n2075), .Q(
        \register[12][23] ) );
  DFFRX1 \register_reg[12][22]  ( .D(n712), .CK(clk), .RN(n2075), .Q(
        \register[12][22] ) );
  DFFRX1 \register_reg[12][21]  ( .D(n711), .CK(clk), .RN(n2075), .Q(
        \register[12][21] ) );
  DFFRX1 \register_reg[12][20]  ( .D(n710), .CK(clk), .RN(n2075), .Q(
        \register[12][20] ) );
  DFFRX1 \register_reg[12][19]  ( .D(n709), .CK(clk), .RN(n2075), .Q(
        \register[12][19] ) );
  DFFRX1 \register_reg[12][18]  ( .D(n708), .CK(clk), .RN(n2075), .Q(
        \register[12][18] ) );
  DFFRX1 \register_reg[12][17]  ( .D(n707), .CK(clk), .RN(n2075), .Q(
        \register[12][17] ) );
  DFFRX1 \register_reg[12][16]  ( .D(n706), .CK(clk), .RN(n2075), .Q(
        \register[12][16] ) );
  DFFRX1 \register_reg[12][15]  ( .D(n705), .CK(clk), .RN(n2074), .Q(
        \register[12][15] ) );
  DFFRX1 \register_reg[12][14]  ( .D(n704), .CK(clk), .RN(n2074), .Q(
        \register[12][14] ) );
  DFFRX1 \register_reg[12][13]  ( .D(n703), .CK(clk), .RN(n2074), .Q(
        \register[12][13] ) );
  DFFRX1 \register_reg[12][12]  ( .D(n702), .CK(clk), .RN(n2074), .Q(
        \register[12][12] ) );
  DFFRX1 \register_reg[12][11]  ( .D(n701), .CK(clk), .RN(n2074), .Q(
        \register[12][11] ) );
  DFFRX1 \register_reg[12][10]  ( .D(n700), .CK(clk), .RN(n2074), .Q(
        \register[12][10] ) );
  DFFRX1 \register_reg[12][9]  ( .D(n699), .CK(clk), .RN(n2074), .Q(
        \register[12][9] ) );
  DFFRX1 \register_reg[16][31]  ( .D(n593), .CK(clk), .RN(n2066), .Q(
        \register[16][31] ) );
  DFFRX1 \register_reg[16][30]  ( .D(n592), .CK(clk), .RN(n2066), .Q(
        \register[16][30] ) );
  DFFRX1 \register_reg[16][29]  ( .D(n591), .CK(clk), .RN(n2066), .Q(
        \register[16][29] ) );
  DFFRX1 \register_reg[16][28]  ( .D(n590), .CK(clk), .RN(n2066), .Q(
        \register[16][28] ) );
  DFFRX1 \register_reg[16][27]  ( .D(n589), .CK(clk), .RN(n2066), .Q(
        \register[16][27] ) );
  DFFRX1 \register_reg[16][26]  ( .D(n588), .CK(clk), .RN(n2065), .Q(
        \register[16][26] ) );
  DFFRX1 \register_reg[16][25]  ( .D(n587), .CK(clk), .RN(n2065), .Q(
        \register[16][25] ) );
  DFFRX1 \register_reg[16][24]  ( .D(n586), .CK(clk), .RN(n2065), .Q(
        \register[16][24] ) );
  DFFRX1 \register_reg[16][23]  ( .D(n585), .CK(clk), .RN(n2065), .Q(
        \register[16][23] ) );
  DFFRX1 \register_reg[16][22]  ( .D(n584), .CK(clk), .RN(n2065), .Q(
        \register[16][22] ) );
  DFFRX1 \register_reg[16][21]  ( .D(n583), .CK(clk), .RN(n2065), .Q(
        \register[16][21] ) );
  DFFRX1 \register_reg[16][20]  ( .D(n582), .CK(clk), .RN(n2065), .Q(
        \register[16][20] ) );
  DFFRX1 \register_reg[16][19]  ( .D(n581), .CK(clk), .RN(n2065), .Q(
        \register[16][19] ) );
  DFFRX1 \register_reg[16][18]  ( .D(n580), .CK(clk), .RN(n2065), .Q(
        \register[16][18] ) );
  DFFRX1 \register_reg[16][17]  ( .D(n579), .CK(clk), .RN(n2065), .Q(
        \register[16][17] ) );
  DFFRX1 \register_reg[16][16]  ( .D(n578), .CK(clk), .RN(n2065), .Q(
        \register[16][16] ) );
  DFFRX1 \register_reg[16][15]  ( .D(n577), .CK(clk), .RN(n2065), .Q(
        \register[16][15] ) );
  DFFRX1 \register_reg[16][14]  ( .D(n576), .CK(clk), .RN(n2065), .Q(
        \register[16][14] ) );
  DFFRX1 \register_reg[16][13]  ( .D(n575), .CK(clk), .RN(n2064), .Q(
        \register[16][13] ) );
  DFFRX1 \register_reg[16][12]  ( .D(n574), .CK(clk), .RN(n2064), .Q(
        \register[16][12] ) );
  DFFRX1 \register_reg[16][11]  ( .D(n573), .CK(clk), .RN(n2064), .Q(
        \register[16][11] ) );
  DFFRX1 \register_reg[16][10]  ( .D(n572), .CK(clk), .RN(n2064), .Q(
        \register[16][10] ) );
  DFFRX1 \register_reg[16][9]  ( .D(n571), .CK(clk), .RN(n2064), .Q(
        \register[16][9] ) );
  DFFRX1 \register_reg[20][31]  ( .D(n465), .CK(clk), .RN(n2056), .Q(
        \register[20][31] ) );
  DFFRX1 \register_reg[20][30]  ( .D(n464), .CK(clk), .RN(n2056), .Q(
        \register[20][30] ) );
  DFFRX1 \register_reg[20][29]  ( .D(n463), .CK(clk), .RN(n2056), .Q(
        \register[20][29] ) );
  DFFRX1 \register_reg[20][28]  ( .D(n462), .CK(clk), .RN(n2056), .Q(
        \register[20][28] ) );
  DFFRX1 \register_reg[20][27]  ( .D(n461), .CK(clk), .RN(n2056), .Q(
        \register[20][27] ) );
  DFFRX1 \register_reg[20][26]  ( .D(n460), .CK(clk), .RN(n2056), .Q(
        \register[20][26] ) );
  DFFRX1 \register_reg[20][25]  ( .D(n459), .CK(clk), .RN(n2056), .Q(
        \register[20][25] ) );
  DFFRX1 \register_reg[20][24]  ( .D(n458), .CK(clk), .RN(n2055), .Q(
        \register[20][24] ) );
  DFFRX1 \register_reg[20][23]  ( .D(n457), .CK(clk), .RN(n2055), .Q(
        \register[20][23] ) );
  DFFRX1 \register_reg[20][22]  ( .D(n456), .CK(clk), .RN(n2055), .Q(
        \register[20][22] ) );
  DFFRX1 \register_reg[20][21]  ( .D(n455), .CK(clk), .RN(n2055), .Q(
        \register[20][21] ) );
  DFFRX1 \register_reg[20][20]  ( .D(n454), .CK(clk), .RN(n2055), .Q(
        \register[20][20] ) );
  DFFRX1 \register_reg[20][19]  ( .D(n453), .CK(clk), .RN(n2055), .Q(
        \register[20][19] ) );
  DFFRX1 \register_reg[20][18]  ( .D(n452), .CK(clk), .RN(n2055), .Q(
        \register[20][18] ) );
  DFFRX1 \register_reg[20][17]  ( .D(n451), .CK(clk), .RN(n2055), .Q(
        \register[20][17] ) );
  DFFRX1 \register_reg[20][16]  ( .D(n450), .CK(clk), .RN(n2055), .Q(
        \register[20][16] ) );
  DFFRX1 \register_reg[20][15]  ( .D(n449), .CK(clk), .RN(n2055), .Q(
        \register[20][15] ) );
  DFFRX1 \register_reg[20][14]  ( .D(n448), .CK(clk), .RN(n2055), .Q(
        \register[20][14] ) );
  DFFRX1 \register_reg[20][13]  ( .D(n447), .CK(clk), .RN(n2055), .Q(
        \register[20][13] ) );
  DFFRX1 \register_reg[20][12]  ( .D(n446), .CK(clk), .RN(n2055), .Q(
        \register[20][12] ) );
  DFFRX1 \register_reg[20][11]  ( .D(n445), .CK(clk), .RN(n2054), .Q(
        \register[20][11] ) );
  DFFRX1 \register_reg[20][10]  ( .D(n444), .CK(clk), .RN(n2054), .Q(
        \register[20][10] ) );
  DFFRX1 \register_reg[20][9]  ( .D(n443), .CK(clk), .RN(n2054), .Q(
        \register[20][9] ) );
  DFFRX1 \register_reg[24][31]  ( .D(n337), .CK(clk), .RN(n2046), .Q(
        \register[24][31] ) );
  DFFRX1 \register_reg[24][30]  ( .D(n336), .CK(clk), .RN(n2046), .Q(
        \register[24][30] ) );
  DFFRX1 \register_reg[24][29]  ( .D(n335), .CK(clk), .RN(n2046), .Q(
        \register[24][29] ) );
  DFFRX1 \register_reg[24][28]  ( .D(n334), .CK(clk), .RN(n2046), .Q(
        \register[24][28] ) );
  DFFRX1 \register_reg[24][27]  ( .D(n333), .CK(clk), .RN(n2046), .Q(
        \register[24][27] ) );
  DFFRX1 \register_reg[24][26]  ( .D(n332), .CK(clk), .RN(n2046), .Q(
        \register[24][26] ) );
  DFFRX1 \register_reg[24][25]  ( .D(n331), .CK(clk), .RN(n2046), .Q(
        \register[24][25] ) );
  DFFRX1 \register_reg[24][24]  ( .D(n330), .CK(clk), .RN(n2046), .Q(
        \register[24][24] ) );
  DFFRX1 \register_reg[24][23]  ( .D(n329), .CK(clk), .RN(n2046), .Q(
        \register[24][23] ) );
  DFFRX1 \register_reg[24][22]  ( .D(n328), .CK(clk), .RN(n2045), .Q(
        \register[24][22] ) );
  DFFRX1 \register_reg[24][21]  ( .D(n327), .CK(clk), .RN(n2045), .Q(
        \register[24][21] ) );
  DFFRX1 \register_reg[24][20]  ( .D(n326), .CK(clk), .RN(n2045), .Q(
        \register[24][20] ) );
  DFFRX1 \register_reg[24][19]  ( .D(n325), .CK(clk), .RN(n2045), .Q(
        \register[24][19] ) );
  DFFRX1 \register_reg[24][18]  ( .D(n324), .CK(clk), .RN(n2045), .Q(
        \register[24][18] ) );
  DFFRX1 \register_reg[24][17]  ( .D(n323), .CK(clk), .RN(n2045), .Q(
        \register[24][17] ) );
  DFFRX1 \register_reg[24][16]  ( .D(n322), .CK(clk), .RN(n2045), .Q(
        \register[24][16] ) );
  DFFRX1 \register_reg[24][15]  ( .D(n321), .CK(clk), .RN(n2045), .Q(
        \register[24][15] ) );
  DFFRX1 \register_reg[24][14]  ( .D(n320), .CK(clk), .RN(n2045), .Q(
        \register[24][14] ) );
  DFFRX1 \register_reg[24][13]  ( .D(n319), .CK(clk), .RN(n2045), .Q(
        \register[24][13] ) );
  DFFRX1 \register_reg[24][12]  ( .D(n318), .CK(clk), .RN(n2045), .Q(
        \register[24][12] ) );
  DFFRX1 \register_reg[24][11]  ( .D(n317), .CK(clk), .RN(n2045), .Q(
        \register[24][11] ) );
  DFFRX1 \register_reg[24][10]  ( .D(n316), .CK(clk), .RN(n2045), .Q(
        \register[24][10] ) );
  DFFRX1 \register_reg[24][9]  ( .D(n315), .CK(clk), .RN(n2044), .Q(
        \register[24][9] ) );
  DFFRX1 \register_reg[28][31]  ( .D(n209), .CK(clk), .RN(n2036), .Q(
        \register[28][31] ) );
  DFFRX1 \register_reg[28][30]  ( .D(n208), .CK(clk), .RN(n2036), .Q(
        \register[28][30] ) );
  DFFRX1 \register_reg[28][29]  ( .D(n207), .CK(clk), .RN(n2036), .Q(
        \register[28][29] ) );
  DFFRX1 \register_reg[28][28]  ( .D(n206), .CK(clk), .RN(n2036), .Q(
        \register[28][28] ) );
  DFFRX1 \register_reg[28][27]  ( .D(n205), .CK(clk), .RN(n2036), .Q(
        \register[28][27] ) );
  DFFRX1 \register_reg[28][26]  ( .D(n204), .CK(clk), .RN(n2036), .Q(
        \register[28][26] ) );
  DFFRX1 \register_reg[28][25]  ( .D(n203), .CK(clk), .RN(n2036), .Q(
        \register[28][25] ) );
  DFFRX1 \register_reg[28][24]  ( .D(n202), .CK(clk), .RN(n2036), .Q(
        \register[28][24] ) );
  DFFRX1 \register_reg[28][23]  ( .D(n201), .CK(clk), .RN(n2036), .Q(
        \register[28][23] ) );
  DFFRX1 \register_reg[28][22]  ( .D(n200), .CK(clk), .RN(n2036), .Q(
        \register[28][22] ) );
  DFFRX1 \register_reg[28][21]  ( .D(n199), .CK(clk), .RN(n2036), .Q(
        \register[28][21] ) );
  DFFRX1 \register_reg[28][20]  ( .D(n198), .CK(clk), .RN(n2035), .Q(
        \register[28][20] ) );
  DFFRX1 \register_reg[28][19]  ( .D(n197), .CK(clk), .RN(n2035), .Q(
        \register[28][19] ) );
  DFFRX1 \register_reg[28][18]  ( .D(n196), .CK(clk), .RN(n2035), .Q(
        \register[28][18] ) );
  DFFRX1 \register_reg[28][17]  ( .D(n195), .CK(clk), .RN(n2035), .Q(
        \register[28][17] ) );
  DFFRX1 \register_reg[28][16]  ( .D(n194), .CK(clk), .RN(n2035), .Q(
        \register[28][16] ) );
  DFFRX1 \register_reg[28][15]  ( .D(n193), .CK(clk), .RN(n2035), .Q(
        \register[28][15] ) );
  DFFRX1 \register_reg[28][14]  ( .D(n192), .CK(clk), .RN(n2035), .Q(
        \register[28][14] ) );
  DFFRX1 \register_reg[28][13]  ( .D(n191), .CK(clk), .RN(n2035), .Q(
        \register[28][13] ) );
  DFFRX1 \register_reg[28][12]  ( .D(n190), .CK(clk), .RN(n2035), .Q(
        \register[28][12] ) );
  DFFRX1 \register_reg[28][11]  ( .D(n189), .CK(clk), .RN(n2035), .Q(
        \register[28][11] ) );
  DFFRX1 \register_reg[28][10]  ( .D(n188), .CK(clk), .RN(n2035), .Q(
        \register[28][10] ) );
  DFFRX1 \register_reg[28][9]  ( .D(n187), .CK(clk), .RN(n2035), .Q(
        \register[28][9] ) );
  DFFRX1 \register_reg[2][31]  ( .D(n1041), .CK(clk), .RN(n2100), .Q(
        \register[2][31] ) );
  DFFRX1 \register_reg[2][30]  ( .D(n1040), .CK(clk), .RN(n2100), .Q(
        \register[2][30] ) );
  DFFRX1 \register_reg[2][29]  ( .D(n1039), .CK(clk), .RN(n2100), .Q(
        \register[2][29] ) );
  DFFRX1 \register_reg[2][28]  ( .D(n1038), .CK(clk), .RN(n2100), .Q(
        \register[2][28] ) );
  DFFRX1 \register_reg[2][27]  ( .D(n1037), .CK(clk), .RN(n2100), .Q(
        \register[2][27] ) );
  DFFRX1 \register_reg[2][26]  ( .D(n1036), .CK(clk), .RN(n2100), .Q(
        \register[2][26] ) );
  DFFRX1 \register_reg[2][25]  ( .D(n1035), .CK(clk), .RN(n2100), .Q(
        \register[2][25] ) );
  DFFRX1 \register_reg[2][24]  ( .D(n1034), .CK(clk), .RN(n2100), .Q(
        \register[2][24] ) );
  DFFRX1 \register_reg[2][23]  ( .D(n1033), .CK(clk), .RN(n2100), .Q(
        \register[2][23] ) );
  DFFRX1 \register_reg[2][22]  ( .D(n1032), .CK(clk), .RN(n2100), .Q(
        \register[2][22] ) );
  DFFRX1 \register_reg[2][21]  ( .D(n1031), .CK(clk), .RN(n2100), .Q(
        \register[2][21] ) );
  DFFRX1 \register_reg[2][20]  ( .D(n1030), .CK(clk), .RN(n2099), .Q(
        \register[2][20] ) );
  DFFRX1 \register_reg[2][19]  ( .D(n1029), .CK(clk), .RN(n2099), .Q(
        \register[2][19] ) );
  DFFRX1 \register_reg[2][18]  ( .D(n1028), .CK(clk), .RN(n2099), .Q(
        \register[2][18] ) );
  DFFRX1 \register_reg[2][17]  ( .D(n1027), .CK(clk), .RN(n2099), .Q(
        \register[2][17] ) );
  DFFRX1 \register_reg[2][16]  ( .D(n1026), .CK(clk), .RN(n2099), .Q(
        \register[2][16] ) );
  DFFRX1 \register_reg[2][15]  ( .D(n1025), .CK(clk), .RN(n2099), .Q(
        \register[2][15] ) );
  DFFRX1 \register_reg[2][14]  ( .D(n1024), .CK(clk), .RN(n2099), .Q(
        \register[2][14] ) );
  DFFRX1 \register_reg[2][13]  ( .D(n1023), .CK(clk), .RN(n2099), .Q(
        \register[2][13] ) );
  DFFRX1 \register_reg[2][12]  ( .D(n1022), .CK(clk), .RN(n2099), .Q(
        \register[2][12] ) );
  DFFRX1 \register_reg[2][11]  ( .D(n1021), .CK(clk), .RN(n2099), .Q(
        \register[2][11] ) );
  DFFRX1 \register_reg[2][10]  ( .D(n1020), .CK(clk), .RN(n2099), .Q(
        \register[2][10] ) );
  DFFRX1 \register_reg[2][9]  ( .D(n1019), .CK(clk), .RN(n2099), .Q(
        \register[2][9] ) );
  DFFRX1 \register_reg[6][31]  ( .D(n913), .CK(clk), .RN(n2090), .Q(
        \register[6][31] ) );
  DFFRX1 \register_reg[6][30]  ( .D(n912), .CK(clk), .RN(n2090), .Q(
        \register[6][30] ) );
  DFFRX1 \register_reg[6][29]  ( .D(n911), .CK(clk), .RN(n2090), .Q(
        \register[6][29] ) );
  DFFRX1 \register_reg[6][28]  ( .D(n910), .CK(clk), .RN(n2090), .Q(
        \register[6][28] ) );
  DFFRX1 \register_reg[6][27]  ( .D(n909), .CK(clk), .RN(n2090), .Q(
        \register[6][27] ) );
  DFFRX1 \register_reg[6][26]  ( .D(n908), .CK(clk), .RN(n2090), .Q(
        \register[6][26] ) );
  DFFRX1 \register_reg[6][25]  ( .D(n907), .CK(clk), .RN(n2090), .Q(
        \register[6][25] ) );
  DFFRX1 \register_reg[6][24]  ( .D(n906), .CK(clk), .RN(n2090), .Q(
        \register[6][24] ) );
  DFFRX1 \register_reg[6][23]  ( .D(n905), .CK(clk), .RN(n2090), .Q(
        \register[6][23] ) );
  DFFRX1 \register_reg[6][22]  ( .D(n904), .CK(clk), .RN(n2090), .Q(
        \register[6][22] ) );
  DFFRX1 \register_reg[6][21]  ( .D(n903), .CK(clk), .RN(n2090), .Q(
        \register[6][21] ) );
  DFFRX1 \register_reg[6][20]  ( .D(n902), .CK(clk), .RN(n2090), .Q(
        \register[6][20] ) );
  DFFRX1 \register_reg[6][19]  ( .D(n901), .CK(clk), .RN(n2090), .Q(
        \register[6][19] ) );
  DFFRX1 \register_reg[6][18]  ( .D(n900), .CK(clk), .RN(n2089), .Q(
        \register[6][18] ) );
  DFFRX1 \register_reg[6][17]  ( .D(n899), .CK(clk), .RN(n2089), .Q(
        \register[6][17] ) );
  DFFRX1 \register_reg[6][16]  ( .D(n898), .CK(clk), .RN(n2089), .Q(
        \register[6][16] ) );
  DFFRX1 \register_reg[6][15]  ( .D(n897), .CK(clk), .RN(n2089), .Q(
        \register[6][15] ) );
  DFFRX1 \register_reg[6][14]  ( .D(n896), .CK(clk), .RN(n2089), .Q(
        \register[6][14] ) );
  DFFRX1 \register_reg[6][13]  ( .D(n895), .CK(clk), .RN(n2089), .Q(
        \register[6][13] ) );
  DFFRX1 \register_reg[6][12]  ( .D(n894), .CK(clk), .RN(n2089), .Q(
        \register[6][12] ) );
  DFFRX1 \register_reg[6][11]  ( .D(n893), .CK(clk), .RN(n2089), .Q(
        \register[6][11] ) );
  DFFRX1 \register_reg[6][10]  ( .D(n892), .CK(clk), .RN(n2089), .Q(
        \register[6][10] ) );
  DFFRX1 \register_reg[6][9]  ( .D(n891), .CK(clk), .RN(n2089), .Q(
        \register[6][9] ) );
  DFFRX1 \register_reg[10][31]  ( .D(n785), .CK(clk), .RN(n2081), .Q(
        \register[10][31] ) );
  DFFRX1 \register_reg[10][30]  ( .D(n784), .CK(clk), .RN(n2081), .Q(
        \register[10][30] ) );
  DFFRX1 \register_reg[10][29]  ( .D(n783), .CK(clk), .RN(n2080), .Q(
        \register[10][29] ) );
  DFFRX1 \register_reg[10][28]  ( .D(n782), .CK(clk), .RN(n2080), .Q(
        \register[10][28] ) );
  DFFRX1 \register_reg[10][27]  ( .D(n781), .CK(clk), .RN(n2080), .Q(
        \register[10][27] ) );
  DFFRX1 \register_reg[10][26]  ( .D(n780), .CK(clk), .RN(n2080), .Q(
        \register[10][26] ) );
  DFFRX1 \register_reg[10][25]  ( .D(n779), .CK(clk), .RN(n2080), .Q(
        \register[10][25] ) );
  DFFRX1 \register_reg[10][24]  ( .D(n778), .CK(clk), .RN(n2080), .Q(
        \register[10][24] ) );
  DFFRX1 \register_reg[10][23]  ( .D(n777), .CK(clk), .RN(n2080), .Q(
        \register[10][23] ) );
  DFFRX1 \register_reg[10][22]  ( .D(n776), .CK(clk), .RN(n2080), .Q(
        \register[10][22] ) );
  DFFRX1 \register_reg[10][21]  ( .D(n775), .CK(clk), .RN(n2080), .Q(
        \register[10][21] ) );
  DFFRX1 \register_reg[10][20]  ( .D(n774), .CK(clk), .RN(n2080), .Q(
        \register[10][20] ) );
  DFFRX1 \register_reg[10][19]  ( .D(n773), .CK(clk), .RN(n2080), .Q(
        \register[10][19] ) );
  DFFRX1 \register_reg[10][18]  ( .D(n772), .CK(clk), .RN(n2080), .Q(
        \register[10][18] ) );
  DFFRX1 \register_reg[10][17]  ( .D(n771), .CK(clk), .RN(n2080), .Q(
        \register[10][17] ) );
  DFFRX1 \register_reg[10][16]  ( .D(n770), .CK(clk), .RN(n2079), .Q(
        \register[10][16] ) );
  DFFRX1 \register_reg[10][15]  ( .D(n769), .CK(clk), .RN(n2079), .Q(
        \register[10][15] ) );
  DFFRX1 \register_reg[10][14]  ( .D(n768), .CK(clk), .RN(n2079), .Q(
        \register[10][14] ) );
  DFFRX1 \register_reg[10][13]  ( .D(n767), .CK(clk), .RN(n2079), .Q(
        \register[10][13] ) );
  DFFRX1 \register_reg[10][12]  ( .D(n766), .CK(clk), .RN(n2079), .Q(
        \register[10][12] ) );
  DFFRX1 \register_reg[10][11]  ( .D(n765), .CK(clk), .RN(n2079), .Q(
        \register[10][11] ) );
  DFFRX1 \register_reg[10][10]  ( .D(n764), .CK(clk), .RN(n2079), .Q(
        \register[10][10] ) );
  DFFRX1 \register_reg[10][9]  ( .D(n763), .CK(clk), .RN(n2079), .Q(
        \register[10][9] ) );
  DFFRX1 \register_reg[14][31]  ( .D(n657), .CK(clk), .RN(n2071), .Q(
        \register[14][31] ) );
  DFFRX1 \register_reg[14][30]  ( .D(n656), .CK(clk), .RN(n2071), .Q(
        \register[14][30] ) );
  DFFRX1 \register_reg[14][29]  ( .D(n655), .CK(clk), .RN(n2071), .Q(
        \register[14][29] ) );
  DFFRX1 \register_reg[14][28]  ( .D(n654), .CK(clk), .RN(n2071), .Q(
        \register[14][28] ) );
  DFFRX1 \register_reg[14][27]  ( .D(n653), .CK(clk), .RN(n2070), .Q(
        \register[14][27] ) );
  DFFRX1 \register_reg[14][26]  ( .D(n652), .CK(clk), .RN(n2070), .Q(
        \register[14][26] ) );
  DFFRX1 \register_reg[14][25]  ( .D(n651), .CK(clk), .RN(n2070), .Q(
        \register[14][25] ) );
  DFFRX1 \register_reg[14][24]  ( .D(n650), .CK(clk), .RN(n2070), .Q(
        \register[14][24] ) );
  DFFRX1 \register_reg[14][23]  ( .D(n649), .CK(clk), .RN(n2070), .Q(
        \register[14][23] ) );
  DFFRX1 \register_reg[14][22]  ( .D(n648), .CK(clk), .RN(n2070), .Q(
        \register[14][22] ) );
  DFFRX1 \register_reg[14][21]  ( .D(n647), .CK(clk), .RN(n2070), .Q(
        \register[14][21] ) );
  DFFRX1 \register_reg[14][20]  ( .D(n646), .CK(clk), .RN(n2070), .Q(
        \register[14][20] ) );
  DFFRX1 \register_reg[14][19]  ( .D(n645), .CK(clk), .RN(n2070), .Q(
        \register[14][19] ) );
  DFFRX1 \register_reg[14][18]  ( .D(n644), .CK(clk), .RN(n2070), .Q(
        \register[14][18] ) );
  DFFRX1 \register_reg[14][17]  ( .D(n643), .CK(clk), .RN(n2070), .Q(
        \register[14][17] ) );
  DFFRX1 \register_reg[14][16]  ( .D(n642), .CK(clk), .RN(n2070), .Q(
        \register[14][16] ) );
  DFFRX1 \register_reg[14][15]  ( .D(n641), .CK(clk), .RN(n2070), .Q(
        \register[14][15] ) );
  DFFRX1 \register_reg[14][14]  ( .D(n640), .CK(clk), .RN(n2069), .Q(
        \register[14][14] ) );
  DFFRX1 \register_reg[14][13]  ( .D(n639), .CK(clk), .RN(n2069), .Q(
        \register[14][13] ) );
  DFFRX1 \register_reg[14][12]  ( .D(n638), .CK(clk), .RN(n2069), .Q(
        \register[14][12] ) );
  DFFRX1 \register_reg[14][11]  ( .D(n637), .CK(clk), .RN(n2069), .Q(
        \register[14][11] ) );
  DFFRX1 \register_reg[14][10]  ( .D(n636), .CK(clk), .RN(n2069), .Q(
        \register[14][10] ) );
  DFFRX1 \register_reg[14][9]  ( .D(n635), .CK(clk), .RN(n2069), .Q(
        \register[14][9] ) );
  DFFRX1 \register_reg[18][31]  ( .D(n529), .CK(clk), .RN(n2061), .Q(
        \register[18][31] ) );
  DFFRX1 \register_reg[18][30]  ( .D(n528), .CK(clk), .RN(n2061), .Q(
        \register[18][30] ) );
  DFFRX1 \register_reg[18][29]  ( .D(n527), .CK(clk), .RN(n2061), .Q(
        \register[18][29] ) );
  DFFRX1 \register_reg[18][28]  ( .D(n526), .CK(clk), .RN(n2061), .Q(
        \register[18][28] ) );
  DFFRX1 \register_reg[18][27]  ( .D(n525), .CK(clk), .RN(n2061), .Q(
        \register[18][27] ) );
  DFFRX1 \register_reg[18][26]  ( .D(n524), .CK(clk), .RN(n2061), .Q(
        \register[18][26] ) );
  DFFRX1 \register_reg[18][25]  ( .D(n523), .CK(clk), .RN(n2060), .Q(
        \register[18][25] ) );
  DFFRX1 \register_reg[18][24]  ( .D(n522), .CK(clk), .RN(n2060), .Q(
        \register[18][24] ) );
  DFFRX1 \register_reg[18][23]  ( .D(n521), .CK(clk), .RN(n2060), .Q(
        \register[18][23] ) );
  DFFRX1 \register_reg[18][22]  ( .D(n520), .CK(clk), .RN(n2060), .Q(
        \register[18][22] ) );
  DFFRX1 \register_reg[18][21]  ( .D(n519), .CK(clk), .RN(n2060), .Q(
        \register[18][21] ) );
  DFFRX1 \register_reg[18][20]  ( .D(n518), .CK(clk), .RN(n2060), .Q(
        \register[18][20] ) );
  DFFRX1 \register_reg[18][19]  ( .D(n517), .CK(clk), .RN(n2060), .Q(
        \register[18][19] ) );
  DFFRX1 \register_reg[18][18]  ( .D(n516), .CK(clk), .RN(n2060), .Q(
        \register[18][18] ) );
  DFFRX1 \register_reg[18][17]  ( .D(n515), .CK(clk), .RN(n2060), .Q(
        \register[18][17] ) );
  DFFRX1 \register_reg[18][16]  ( .D(n514), .CK(clk), .RN(n2060), .Q(
        \register[18][16] ) );
  DFFRX1 \register_reg[18][15]  ( .D(n513), .CK(clk), .RN(n2060), .Q(
        \register[18][15] ) );
  DFFRX1 \register_reg[18][14]  ( .D(n512), .CK(clk), .RN(n2060), .Q(
        \register[18][14] ) );
  DFFRX1 \register_reg[18][13]  ( .D(n511), .CK(clk), .RN(n2060), .Q(
        \register[18][13] ) );
  DFFRX1 \register_reg[18][12]  ( .D(n510), .CK(clk), .RN(n2059), .Q(
        \register[18][12] ) );
  DFFRX1 \register_reg[18][11]  ( .D(n509), .CK(clk), .RN(n2059), .Q(
        \register[18][11] ) );
  DFFRX1 \register_reg[18][10]  ( .D(n508), .CK(clk), .RN(n2059), .Q(
        \register[18][10] ) );
  DFFRX1 \register_reg[18][9]  ( .D(n507), .CK(clk), .RN(n2059), .Q(
        \register[18][9] ) );
  DFFRX1 \register_reg[22][31]  ( .D(n401), .CK(clk), .RN(n2051), .Q(
        \register[22][31] ) );
  DFFRX1 \register_reg[22][30]  ( .D(n400), .CK(clk), .RN(n2051), .Q(
        \register[22][30] ) );
  DFFRX1 \register_reg[22][29]  ( .D(n399), .CK(clk), .RN(n2051), .Q(
        \register[22][29] ) );
  DFFRX1 \register_reg[22][28]  ( .D(n398), .CK(clk), .RN(n2051), .Q(
        \register[22][28] ) );
  DFFRX1 \register_reg[22][27]  ( .D(n397), .CK(clk), .RN(n2051), .Q(
        \register[22][27] ) );
  DFFRX1 \register_reg[22][26]  ( .D(n396), .CK(clk), .RN(n2051), .Q(
        \register[22][26] ) );
  DFFRX1 \register_reg[22][25]  ( .D(n395), .CK(clk), .RN(n2051), .Q(
        \register[22][25] ) );
  DFFRX1 \register_reg[22][24]  ( .D(n394), .CK(clk), .RN(n2051), .Q(
        \register[22][24] ) );
  DFFRX1 \register_reg[22][23]  ( .D(n393), .CK(clk), .RN(n2050), .Q(
        \register[22][23] ) );
  DFFRX1 \register_reg[22][22]  ( .D(n392), .CK(clk), .RN(n2050), .Q(
        \register[22][22] ) );
  DFFRX1 \register_reg[22][21]  ( .D(n391), .CK(clk), .RN(n2050), .Q(
        \register[22][21] ) );
  DFFRX1 \register_reg[22][20]  ( .D(n390), .CK(clk), .RN(n2050), .Q(
        \register[22][20] ) );
  DFFRX1 \register_reg[22][19]  ( .D(n389), .CK(clk), .RN(n2050), .Q(
        \register[22][19] ) );
  DFFRX1 \register_reg[22][18]  ( .D(n388), .CK(clk), .RN(n2050), .Q(
        \register[22][18] ) );
  DFFRX1 \register_reg[22][17]  ( .D(n387), .CK(clk), .RN(n2050), .Q(
        \register[22][17] ) );
  DFFRX1 \register_reg[22][16]  ( .D(n386), .CK(clk), .RN(n2050), .Q(
        \register[22][16] ) );
  DFFRX1 \register_reg[22][15]  ( .D(n385), .CK(clk), .RN(n2050), .Q(
        \register[22][15] ) );
  DFFRX1 \register_reg[22][14]  ( .D(n384), .CK(clk), .RN(n2050), .Q(
        \register[22][14] ) );
  DFFRX1 \register_reg[22][13]  ( .D(n383), .CK(clk), .RN(n2050), .Q(
        \register[22][13] ) );
  DFFRX1 \register_reg[22][12]  ( .D(n382), .CK(clk), .RN(n2050), .Q(
        \register[22][12] ) );
  DFFRX1 \register_reg[22][11]  ( .D(n381), .CK(clk), .RN(n2050), .Q(
        \register[22][11] ) );
  DFFRX1 \register_reg[22][10]  ( .D(n380), .CK(clk), .RN(n2049), .Q(
        \register[22][10] ) );
  DFFRX1 \register_reg[22][9]  ( .D(n379), .CK(clk), .RN(n2049), .Q(
        \register[22][9] ) );
  DFFRX1 \register_reg[26][31]  ( .D(n273), .CK(clk), .RN(n2041), .Q(
        \register[26][31] ) );
  DFFRX1 \register_reg[26][30]  ( .D(n272), .CK(clk), .RN(n2041), .Q(
        \register[26][30] ) );
  DFFRX1 \register_reg[26][29]  ( .D(n271), .CK(clk), .RN(n2041), .Q(
        \register[26][29] ) );
  DFFRX1 \register_reg[26][28]  ( .D(n270), .CK(clk), .RN(n2041), .Q(
        \register[26][28] ) );
  DFFRX1 \register_reg[26][27]  ( .D(n269), .CK(clk), .RN(n2041), .Q(
        \register[26][27] ) );
  DFFRX1 \register_reg[26][26]  ( .D(n268), .CK(clk), .RN(n2041), .Q(
        \register[26][26] ) );
  DFFRX1 \register_reg[26][25]  ( .D(n267), .CK(clk), .RN(n2041), .Q(
        \register[26][25] ) );
  DFFRX1 \register_reg[26][24]  ( .D(n266), .CK(clk), .RN(n2041), .Q(
        \register[26][24] ) );
  DFFRX1 \register_reg[26][23]  ( .D(n265), .CK(clk), .RN(n2041), .Q(
        \register[26][23] ) );
  DFFRX1 \register_reg[26][22]  ( .D(n264), .CK(clk), .RN(n2041), .Q(
        \register[26][22] ) );
  DFFRX1 \register_reg[26][21]  ( .D(n263), .CK(clk), .RN(n2040), .Q(
        \register[26][21] ) );
  DFFRX1 \register_reg[26][20]  ( .D(n262), .CK(clk), .RN(n2040), .Q(
        \register[26][20] ) );
  DFFRX1 \register_reg[26][19]  ( .D(n261), .CK(clk), .RN(n2040), .Q(
        \register[26][19] ) );
  DFFRX1 \register_reg[26][18]  ( .D(n260), .CK(clk), .RN(n2040), .Q(
        \register[26][18] ) );
  DFFRX1 \register_reg[26][17]  ( .D(n259), .CK(clk), .RN(n2040), .Q(
        \register[26][17] ) );
  DFFRX1 \register_reg[26][16]  ( .D(n258), .CK(clk), .RN(n2040), .Q(
        \register[26][16] ) );
  DFFRX1 \register_reg[26][15]  ( .D(n257), .CK(clk), .RN(n2040), .Q(
        \register[26][15] ) );
  DFFRX1 \register_reg[26][14]  ( .D(n256), .CK(clk), .RN(n2040), .Q(
        \register[26][14] ) );
  DFFRX1 \register_reg[26][13]  ( .D(n255), .CK(clk), .RN(n2040), .Q(
        \register[26][13] ) );
  DFFRX1 \register_reg[26][12]  ( .D(n254), .CK(clk), .RN(n2040), .Q(
        \register[26][12] ) );
  DFFRX1 \register_reg[26][11]  ( .D(n253), .CK(clk), .RN(n2040), .Q(
        \register[26][11] ) );
  DFFRX1 \register_reg[26][10]  ( .D(n252), .CK(clk), .RN(n2040), .Q(
        \register[26][10] ) );
  DFFRX1 \register_reg[26][9]  ( .D(n251), .CK(clk), .RN(n2040), .Q(
        \register[26][9] ) );
  DFFRX1 \register_reg[30][31]  ( .D(n145), .CK(clk), .RN(n2031), .Q(
        \register[30][31] ) );
  DFFRX1 \register_reg[30][30]  ( .D(n144), .CK(clk), .RN(n2031), .Q(
        \register[30][30] ) );
  DFFRX1 \register_reg[30][29]  ( .D(n143), .CK(clk), .RN(n2031), .Q(
        \register[30][29] ) );
  DFFRX1 \register_reg[30][28]  ( .D(n142), .CK(clk), .RN(n2031), .Q(
        \register[30][28] ) );
  DFFRX1 \register_reg[30][27]  ( .D(n141), .CK(clk), .RN(n2031), .Q(
        \register[30][27] ) );
  DFFRX1 \register_reg[30][26]  ( .D(n140), .CK(clk), .RN(n2031), .Q(
        \register[30][26] ) );
  DFFRX1 \register_reg[30][25]  ( .D(n139), .CK(clk), .RN(n2031), .Q(
        \register[30][25] ) );
  DFFRX1 \register_reg[30][24]  ( .D(n138), .CK(clk), .RN(n2031), .Q(
        \register[30][24] ) );
  DFFRX1 \register_reg[30][23]  ( .D(n137), .CK(clk), .RN(n2031), .Q(
        \register[30][23] ) );
  DFFRX1 \register_reg[30][22]  ( .D(n136), .CK(clk), .RN(n2031), .Q(
        \register[30][22] ) );
  DFFRX1 \register_reg[30][21]  ( .D(n135), .CK(clk), .RN(n2031), .Q(
        \register[30][21] ) );
  DFFRX1 \register_reg[30][20]  ( .D(n134), .CK(clk), .RN(n2031), .Q(
        \register[30][20] ) );
  DFFRX1 \register_reg[30][19]  ( .D(n133), .CK(clk), .RN(n2030), .Q(
        \register[30][19] ) );
  DFFRX1 \register_reg[30][18]  ( .D(n132), .CK(clk), .RN(n2030), .Q(
        \register[30][18] ) );
  DFFRX1 \register_reg[30][17]  ( .D(n131), .CK(clk), .RN(n2030), .Q(
        \register[30][17] ) );
  DFFRX1 \register_reg[30][16]  ( .D(n130), .CK(clk), .RN(n2030), .Q(
        \register[30][16] ) );
  DFFRX1 \register_reg[30][15]  ( .D(n129), .CK(clk), .RN(n2030), .Q(
        \register[30][15] ) );
  DFFRX1 \register_reg[30][14]  ( .D(n128), .CK(clk), .RN(n2030), .Q(
        \register[30][14] ) );
  DFFRX1 \register_reg[30][13]  ( .D(n127), .CK(clk), .RN(n2030), .Q(
        \register[30][13] ) );
  DFFRX1 \register_reg[30][12]  ( .D(n126), .CK(clk), .RN(n2030), .Q(
        \register[30][12] ) );
  DFFRX1 \register_reg[30][11]  ( .D(n125), .CK(clk), .RN(n2030), .Q(
        \register[30][11] ) );
  DFFRX1 \register_reg[30][10]  ( .D(n124), .CK(clk), .RN(n2030), .Q(
        \register[30][10] ) );
  DFFRX1 \register_reg[30][9]  ( .D(n123), .CK(clk), .RN(n2030), .Q(
        \register[30][9] ) );
  DFFRX1 \register_reg[3][8]  ( .D(n986), .CK(clk), .RN(n2096), .Q(
        \register[3][8] ) );
  DFFRX1 \register_reg[3][7]  ( .D(n985), .CK(clk), .RN(n2096), .Q(
        \register[3][7] ) );
  DFFRX1 \register_reg[3][6]  ( .D(n984), .CK(clk), .RN(n2096), .Q(
        \register[3][6] ) );
  DFFRX1 \register_reg[3][5]  ( .D(n983), .CK(clk), .RN(n2096), .Q(
        \register[3][5] ) );
  DFFRX1 \register_reg[3][4]  ( .D(n982), .CK(clk), .RN(n2096), .Q(
        \register[3][4] ) );
  DFFRX1 \register_reg[7][8]  ( .D(n858), .CK(clk), .RN(n2086), .Q(
        \register[7][8] ) );
  DFFRX1 \register_reg[7][7]  ( .D(n857), .CK(clk), .RN(n2086), .Q(
        \register[7][7] ) );
  DFFRX1 \register_reg[7][6]  ( .D(n856), .CK(clk), .RN(n2086), .Q(
        \register[7][6] ) );
  DFFRX1 \register_reg[7][5]  ( .D(n855), .CK(clk), .RN(n2086), .Q(
        \register[7][5] ) );
  DFFRX1 \register_reg[7][4]  ( .D(n854), .CK(clk), .RN(n2086), .Q(
        \register[7][4] ) );
  DFFRX1 \register_reg[11][8]  ( .D(n730), .CK(clk), .RN(n2076), .Q(
        \register[11][8] ) );
  DFFRX1 \register_reg[11][7]  ( .D(n729), .CK(clk), .RN(n2076), .Q(
        \register[11][7] ) );
  DFFRX1 \register_reg[11][6]  ( .D(n728), .CK(clk), .RN(n2076), .Q(
        \register[11][6] ) );
  DFFRX1 \register_reg[11][5]  ( .D(n727), .CK(clk), .RN(n2076), .Q(
        \register[11][5] ) );
  DFFRX1 \register_reg[11][4]  ( .D(n726), .CK(clk), .RN(n2076), .Q(
        \register[11][4] ) );
  DFFRX1 \register_reg[15][8]  ( .D(n602), .CK(clk), .RN(n2067), .Q(
        \register[15][8] ) );
  DFFRX1 \register_reg[15][7]  ( .D(n601), .CK(clk), .RN(n2066), .Q(
        \register[15][7] ) );
  DFFRX1 \register_reg[15][6]  ( .D(n600), .CK(clk), .RN(n2066), .Q(
        \register[15][6] ) );
  DFFRX1 \register_reg[15][5]  ( .D(n599), .CK(clk), .RN(n2066), .Q(
        \register[15][5] ) );
  DFFRX1 \register_reg[15][4]  ( .D(n598), .CK(clk), .RN(n2066), .Q(
        \register[15][4] ) );
  DFFRX1 \register_reg[19][8]  ( .D(n474), .CK(clk), .RN(n2057), .Q(
        \register[19][8] ) );
  DFFRX1 \register_reg[19][7]  ( .D(n473), .CK(clk), .RN(n2057), .Q(
        \register[19][7] ) );
  DFFRX1 \register_reg[19][6]  ( .D(n472), .CK(clk), .RN(n2057), .Q(
        \register[19][6] ) );
  DFFRX1 \register_reg[19][5]  ( .D(n471), .CK(clk), .RN(n2056), .Q(
        \register[19][5] ) );
  DFFRX1 \register_reg[19][4]  ( .D(n470), .CK(clk), .RN(n2056), .Q(
        \register[19][4] ) );
  DFFRX1 \register_reg[23][8]  ( .D(n346), .CK(clk), .RN(n2047), .Q(
        \register[23][8] ) );
  DFFRX1 \register_reg[23][7]  ( .D(n345), .CK(clk), .RN(n2047), .Q(
        \register[23][7] ) );
  DFFRX1 \register_reg[23][6]  ( .D(n344), .CK(clk), .RN(n2047), .Q(
        \register[23][6] ) );
  DFFRX1 \register_reg[23][5]  ( .D(n343), .CK(clk), .RN(n2047), .Q(
        \register[23][5] ) );
  DFFRX1 \register_reg[23][4]  ( .D(n342), .CK(clk), .RN(n2047), .Q(
        \register[23][4] ) );
  DFFRX1 \register_reg[31][8]  ( .D(n90), .CK(clk), .RN(n2027), .Q(
        \register[31][8] ) );
  DFFRX1 \register_reg[31][7]  ( .D(n89), .CK(clk), .RN(n2027), .Q(
        \register[31][7] ) );
  DFFRX1 \register_reg[31][6]  ( .D(n88), .CK(clk), .RN(n2027), .Q(
        \register[31][6] ) );
  DFFRX1 \register_reg[31][5]  ( .D(n87), .CK(clk), .RN(n2027), .Q(
        \register[31][5] ) );
  DFFRX1 \register_reg[31][4]  ( .D(n86), .CK(clk), .RN(n2027), .Q(
        \register[31][4] ) );
  DFFRX1 \register_reg[1][8]  ( .D(n1050), .CK(clk), .RN(n2101), .Q(
        \register[1][8] ) );
  DFFRX1 \register_reg[1][7]  ( .D(n1049), .CK(clk), .RN(n2101), .Q(
        \register[1][7] ) );
  DFFRX1 \register_reg[1][6]  ( .D(n1048), .CK(clk), .RN(n2101), .Q(
        \register[1][6] ) );
  DFFRX1 \register_reg[1][5]  ( .D(n1047), .CK(clk), .RN(n2101), .Q(
        \register[1][5] ) );
  DFFRX1 \register_reg[1][4]  ( .D(n1046), .CK(clk), .RN(n2101), .Q(
        \register[1][4] ) );
  DFFRX1 \register_reg[5][8]  ( .D(n922), .CK(clk), .RN(n2091), .Q(
        \register[5][8] ) );
  DFFRX1 \register_reg[5][7]  ( .D(n921), .CK(clk), .RN(n2091), .Q(
        \register[5][7] ) );
  DFFRX1 \register_reg[5][6]  ( .D(n920), .CK(clk), .RN(n2091), .Q(
        \register[5][6] ) );
  DFFRX1 \register_reg[5][5]  ( .D(n919), .CK(clk), .RN(n2091), .Q(
        \register[5][5] ) );
  DFFRX1 \register_reg[5][4]  ( .D(n918), .CK(clk), .RN(n2091), .Q(
        \register[5][4] ) );
  DFFRX1 \register_reg[9][8]  ( .D(n794), .CK(clk), .RN(n2081), .Q(
        \register[9][8] ) );
  DFFRX1 \register_reg[9][7]  ( .D(n793), .CK(clk), .RN(n2081), .Q(
        \register[9][7] ) );
  DFFRX1 \register_reg[9][6]  ( .D(n792), .CK(clk), .RN(n2081), .Q(
        \register[9][6] ) );
  DFFRX1 \register_reg[9][5]  ( .D(n791), .CK(clk), .RN(n2081), .Q(
        \register[9][5] ) );
  DFFRX1 \register_reg[9][4]  ( .D(n790), .CK(clk), .RN(n2081), .Q(
        \register[9][4] ) );
  DFFRX1 \register_reg[13][8]  ( .D(n666), .CK(clk), .RN(n2071), .Q(
        \register[13][8] ) );
  DFFRX1 \register_reg[13][7]  ( .D(n665), .CK(clk), .RN(n2071), .Q(
        \register[13][7] ) );
  DFFRX1 \register_reg[13][6]  ( .D(n664), .CK(clk), .RN(n2071), .Q(
        \register[13][6] ) );
  DFFRX1 \register_reg[13][5]  ( .D(n663), .CK(clk), .RN(n2071), .Q(
        \register[13][5] ) );
  DFFRX1 \register_reg[13][4]  ( .D(n662), .CK(clk), .RN(n2071), .Q(
        \register[13][4] ) );
  DFFRX1 \register_reg[17][8]  ( .D(n538), .CK(clk), .RN(n2062), .Q(
        \register[17][8] ) );
  DFFRX1 \register_reg[17][7]  ( .D(n537), .CK(clk), .RN(n2062), .Q(
        \register[17][7] ) );
  DFFRX1 \register_reg[17][6]  ( .D(n536), .CK(clk), .RN(n2061), .Q(
        \register[17][6] ) );
  DFFRX1 \register_reg[17][5]  ( .D(n535), .CK(clk), .RN(n2061), .Q(
        \register[17][5] ) );
  DFFRX1 \register_reg[17][4]  ( .D(n534), .CK(clk), .RN(n2061), .Q(
        \register[17][4] ) );
  DFFRX1 \register_reg[21][8]  ( .D(n410), .CK(clk), .RN(n2052), .Q(
        \register[21][8] ) );
  DFFRX1 \register_reg[21][7]  ( .D(n409), .CK(clk), .RN(n2052), .Q(
        \register[21][7] ) );
  DFFRX1 \register_reg[21][6]  ( .D(n408), .CK(clk), .RN(n2052), .Q(
        \register[21][6] ) );
  DFFRX1 \register_reg[21][5]  ( .D(n407), .CK(clk), .RN(n2052), .Q(
        \register[21][5] ) );
  DFFRX1 \register_reg[21][4]  ( .D(n406), .CK(clk), .RN(n2051), .Q(
        \register[21][4] ) );
  DFFRX1 \register_reg[0][8]  ( .D(n1082), .CK(clk), .RN(n2103), .Q(
        \register[0][8] ) );
  DFFRX1 \register_reg[0][7]  ( .D(n1081), .CK(clk), .RN(n2103), .Q(
        \register[0][7] ) );
  DFFRX1 \register_reg[0][6]  ( .D(n1080), .CK(clk), .RN(n2103), .Q(
        \register[0][6] ) );
  DFFRX1 \register_reg[0][5]  ( .D(n1079), .CK(clk), .RN(n2103), .Q(
        \register[0][5] ) );
  DFFRX1 \register_reg[0][4]  ( .D(n1078), .CK(clk), .RN(n2103), .Q(
        \register[0][4] ) );
  DFFRX1 \register_reg[4][8]  ( .D(n954), .CK(clk), .RN(n2094), .Q(
        \register[4][8] ) );
  DFFRX1 \register_reg[4][7]  ( .D(n953), .CK(clk), .RN(n2094), .Q(
        \register[4][7] ) );
  DFFRX1 \register_reg[4][6]  ( .D(n952), .CK(clk), .RN(n2093), .Q(
        \register[4][6] ) );
  DFFRX1 \register_reg[4][5]  ( .D(n951), .CK(clk), .RN(n2093), .Q(
        \register[4][5] ) );
  DFFRX1 \register_reg[4][4]  ( .D(n950), .CK(clk), .RN(n2093), .Q(
        \register[4][4] ) );
  DFFRX1 \register_reg[8][8]  ( .D(n826), .CK(clk), .RN(n2084), .Q(
        \register[8][8] ) );
  DFFRX1 \register_reg[8][7]  ( .D(n825), .CK(clk), .RN(n2084), .Q(
        \register[8][7] ) );
  DFFRX1 \register_reg[8][6]  ( .D(n824), .CK(clk), .RN(n2084), .Q(
        \register[8][6] ) );
  DFFRX1 \register_reg[8][5]  ( .D(n823), .CK(clk), .RN(n2084), .Q(
        \register[8][5] ) );
  DFFRX1 \register_reg[8][4]  ( .D(n822), .CK(clk), .RN(n2083), .Q(
        \register[8][4] ) );
  DFFRX1 \register_reg[12][8]  ( .D(n698), .CK(clk), .RN(n2074), .Q(
        \register[12][8] ) );
  DFFRX1 \register_reg[12][7]  ( .D(n697), .CK(clk), .RN(n2074), .Q(
        \register[12][7] ) );
  DFFRX1 \register_reg[12][6]  ( .D(n696), .CK(clk), .RN(n2074), .Q(
        \register[12][6] ) );
  DFFRX1 \register_reg[12][5]  ( .D(n695), .CK(clk), .RN(n2074), .Q(
        \register[12][5] ) );
  DFFRX1 \register_reg[12][4]  ( .D(n694), .CK(clk), .RN(n2074), .Q(
        \register[12][4] ) );
  DFFRX1 \register_reg[16][8]  ( .D(n570), .CK(clk), .RN(n2064), .Q(
        \register[16][8] ) );
  DFFRX1 \register_reg[16][7]  ( .D(n569), .CK(clk), .RN(n2064), .Q(
        \register[16][7] ) );
  DFFRX1 \register_reg[16][6]  ( .D(n568), .CK(clk), .RN(n2064), .Q(
        \register[16][6] ) );
  DFFRX1 \register_reg[16][5]  ( .D(n567), .CK(clk), .RN(n2064), .Q(
        \register[16][5] ) );
  DFFRX1 \register_reg[16][4]  ( .D(n566), .CK(clk), .RN(n2064), .Q(
        \register[16][4] ) );
  DFFRX1 \register_reg[20][8]  ( .D(n442), .CK(clk), .RN(n2054), .Q(
        \register[20][8] ) );
  DFFRX1 \register_reg[20][7]  ( .D(n441), .CK(clk), .RN(n2054), .Q(
        \register[20][7] ) );
  DFFRX1 \register_reg[20][6]  ( .D(n440), .CK(clk), .RN(n2054), .Q(
        \register[20][6] ) );
  DFFRX1 \register_reg[20][5]  ( .D(n439), .CK(clk), .RN(n2054), .Q(
        \register[20][5] ) );
  DFFRX1 \register_reg[20][4]  ( .D(n438), .CK(clk), .RN(n2054), .Q(
        \register[20][4] ) );
  DFFRX1 \register_reg[24][5]  ( .D(n311), .CK(clk), .RN(n2044), .Q(
        \register[24][5] ) );
  DFFRX1 \register_reg[24][4]  ( .D(n310), .CK(clk), .RN(n2044), .Q(
        \register[24][4] ) );
  DFFRX1 \register_reg[2][8]  ( .D(n1018), .CK(clk), .RN(n2099), .Q(
        \register[2][8] ) );
  DFFRX1 \register_reg[2][7]  ( .D(n1017), .CK(clk), .RN(n2098), .Q(
        \register[2][7] ) );
  DFFRX1 \register_reg[2][6]  ( .D(n1016), .CK(clk), .RN(n2098), .Q(
        \register[2][6] ) );
  DFFRX1 \register_reg[2][5]  ( .D(n1015), .CK(clk), .RN(n2098), .Q(
        \register[2][5] ) );
  DFFRX1 \register_reg[2][4]  ( .D(n1014), .CK(clk), .RN(n2098), .Q(
        \register[2][4] ) );
  DFFRX1 \register_reg[6][8]  ( .D(n890), .CK(clk), .RN(n2089), .Q(
        \register[6][8] ) );
  DFFRX1 \register_reg[6][7]  ( .D(n889), .CK(clk), .RN(n2089), .Q(
        \register[6][7] ) );
  DFFRX1 \register_reg[6][6]  ( .D(n888), .CK(clk), .RN(n2089), .Q(
        \register[6][6] ) );
  DFFRX1 \register_reg[6][5]  ( .D(n887), .CK(clk), .RN(n2088), .Q(
        \register[6][5] ) );
  DFFRX1 \register_reg[6][4]  ( .D(n886), .CK(clk), .RN(n2088), .Q(
        \register[6][4] ) );
  DFFRX1 \register_reg[10][8]  ( .D(n762), .CK(clk), .RN(n2079), .Q(
        \register[10][8] ) );
  DFFRX1 \register_reg[10][7]  ( .D(n761), .CK(clk), .RN(n2079), .Q(
        \register[10][7] ) );
  DFFRX1 \register_reg[10][6]  ( .D(n760), .CK(clk), .RN(n2079), .Q(
        \register[10][6] ) );
  DFFRX1 \register_reg[10][5]  ( .D(n759), .CK(clk), .RN(n2079), .Q(
        \register[10][5] ) );
  DFFRX1 \register_reg[10][4]  ( .D(n758), .CK(clk), .RN(n2079), .Q(
        \register[10][4] ) );
  DFFRX1 \register_reg[14][8]  ( .D(n634), .CK(clk), .RN(n2069), .Q(
        \register[14][8] ) );
  DFFRX1 \register_reg[14][7]  ( .D(n633), .CK(clk), .RN(n2069), .Q(
        \register[14][7] ) );
  DFFRX1 \register_reg[14][6]  ( .D(n632), .CK(clk), .RN(n2069), .Q(
        \register[14][6] ) );
  DFFRX1 \register_reg[14][5]  ( .D(n631), .CK(clk), .RN(n2069), .Q(
        \register[14][5] ) );
  DFFRX1 \register_reg[14][4]  ( .D(n630), .CK(clk), .RN(n2069), .Q(
        \register[14][4] ) );
  DFFRX1 \register_reg[18][8]  ( .D(n506), .CK(clk), .RN(n2059), .Q(
        \register[18][8] ) );
  DFFRX1 \register_reg[18][7]  ( .D(n505), .CK(clk), .RN(n2059), .Q(
        \register[18][7] ) );
  DFFRX1 \register_reg[18][6]  ( .D(n504), .CK(clk), .RN(n2059), .Q(
        \register[18][6] ) );
  DFFRX1 \register_reg[18][5]  ( .D(n503), .CK(clk), .RN(n2059), .Q(
        \register[18][5] ) );
  DFFRX1 \register_reg[18][4]  ( .D(n502), .CK(clk), .RN(n2059), .Q(
        \register[18][4] ) );
  DFFRX1 \register_reg[22][8]  ( .D(n378), .CK(clk), .RN(n2049), .Q(
        \register[22][8] ) );
  DFFRX1 \register_reg[22][7]  ( .D(n377), .CK(clk), .RN(n2049), .Q(
        \register[22][7] ) );
  DFFRX1 \register_reg[22][6]  ( .D(n376), .CK(clk), .RN(n2049), .Q(
        \register[22][6] ) );
  DFFRX1 \register_reg[22][5]  ( .D(n375), .CK(clk), .RN(n2049), .Q(
        \register[22][5] ) );
  DFFRX1 \register_reg[22][4]  ( .D(n374), .CK(clk), .RN(n2049), .Q(
        \register[22][4] ) );
  DFFRX1 \register_reg[3][3]  ( .D(n981), .CK(clk), .RN(n2096), .Q(
        \register[3][3] ) );
  DFFRX1 \register_reg[3][2]  ( .D(n980), .CK(clk), .RN(n2096), .Q(
        \register[3][2] ) );
  DFFRX1 \register_reg[3][1]  ( .D(n979), .CK(clk), .RN(n2096), .Q(
        \register[3][1] ) );
  DFFRX1 \register_reg[3][0]  ( .D(n978), .CK(clk), .RN(n2095), .Q(
        \register[3][0] ) );
  DFFRX1 \register_reg[7][3]  ( .D(n853), .CK(clk), .RN(n2086), .Q(
        \register[7][3] ) );
  DFFRX1 \register_reg[7][2]  ( .D(n852), .CK(clk), .RN(n2086), .Q(
        \register[7][2] ) );
  DFFRX1 \register_reg[7][1]  ( .D(n851), .CK(clk), .RN(n2086), .Q(
        \register[7][1] ) );
  DFFRX1 \register_reg[7][0]  ( .D(n850), .CK(clk), .RN(n2086), .Q(
        \register[7][0] ) );
  DFFRX1 \register_reg[11][3]  ( .D(n725), .CK(clk), .RN(n2076), .Q(
        \register[11][3] ) );
  DFFRX1 \register_reg[11][2]  ( .D(n724), .CK(clk), .RN(n2076), .Q(
        \register[11][2] ) );
  DFFRX1 \register_reg[11][1]  ( .D(n723), .CK(clk), .RN(n2076), .Q(
        \register[11][1] ) );
  DFFRX1 \register_reg[11][0]  ( .D(n722), .CK(clk), .RN(n2076), .Q(
        \register[11][0] ) );
  DFFRX1 \register_reg[15][3]  ( .D(n597), .CK(clk), .RN(n2066), .Q(
        \register[15][3] ) );
  DFFRX1 \register_reg[15][2]  ( .D(n596), .CK(clk), .RN(n2066), .Q(
        \register[15][2] ) );
  DFFRX1 \register_reg[15][1]  ( .D(n595), .CK(clk), .RN(n2066), .Q(
        \register[15][1] ) );
  DFFRX1 \register_reg[15][0]  ( .D(n594), .CK(clk), .RN(n2066), .Q(
        \register[15][0] ) );
  DFFRX1 \register_reg[19][3]  ( .D(n469), .CK(clk), .RN(n2056), .Q(
        \register[19][3] ) );
  DFFRX1 \register_reg[19][2]  ( .D(n468), .CK(clk), .RN(n2056), .Q(
        \register[19][2] ) );
  DFFRX1 \register_reg[19][1]  ( .D(n467), .CK(clk), .RN(n2056), .Q(
        \register[19][1] ) );
  DFFRX1 \register_reg[19][0]  ( .D(n466), .CK(clk), .RN(n2056), .Q(
        \register[19][0] ) );
  DFFRX1 \register_reg[23][3]  ( .D(n341), .CK(clk), .RN(n2046), .Q(
        \register[23][3] ) );
  DFFRX1 \register_reg[23][2]  ( .D(n340), .CK(clk), .RN(n2046), .Q(
        \register[23][2] ) );
  DFFRX1 \register_reg[23][1]  ( .D(n339), .CK(clk), .RN(n2046), .Q(
        \register[23][1] ) );
  DFFRX1 \register_reg[23][0]  ( .D(n338), .CK(clk), .RN(n2046), .Q(
        \register[23][0] ) );
  DFFRX1 \register_reg[27][2]  ( .D(n212), .CK(clk), .RN(n2037), .Q(
        \register[27][2] ) );
  DFFRX1 \register_reg[27][1]  ( .D(n211), .CK(clk), .RN(n2036), .Q(
        \register[27][1] ) );
  DFFRX1 \register_reg[27][0]  ( .D(n210), .CK(clk), .RN(n2036), .Q(
        \register[27][0] ) );
  DFFRX1 \register_reg[31][3]  ( .D(n85), .CK(clk), .RN(n2027), .Q(
        \register[31][3] ) );
  DFFRX1 \register_reg[31][2]  ( .D(n84), .CK(clk), .RN(n2027), .Q(
        \register[31][2] ) );
  DFFRX1 \register_reg[31][1]  ( .D(n83), .CK(clk), .RN(n2027), .Q(
        \register[31][1] ) );
  DFFRX1 \register_reg[31][0]  ( .D(n82), .CK(clk), .RN(n2027), .Q(
        \register[31][0] ) );
  DFFRX1 \register_reg[1][3]  ( .D(n1045), .CK(clk), .RN(n2101), .Q(
        \register[1][3] ) );
  DFFRX1 \register_reg[1][2]  ( .D(n1044), .CK(clk), .RN(n2101), .Q(
        \register[1][2] ) );
  DFFRX1 \register_reg[1][1]  ( .D(n1043), .CK(clk), .RN(n2100), .Q(
        \register[1][1] ) );
  DFFRX1 \register_reg[1][0]  ( .D(n1042), .CK(clk), .RN(n2100), .Q(
        \register[1][0] ) );
  DFFRX1 \register_reg[5][3]  ( .D(n917), .CK(clk), .RN(n2091), .Q(
        \register[5][3] ) );
  DFFRX1 \register_reg[5][2]  ( .D(n916), .CK(clk), .RN(n2091), .Q(
        \register[5][2] ) );
  DFFRX1 \register_reg[5][1]  ( .D(n915), .CK(clk), .RN(n2091), .Q(
        \register[5][1] ) );
  DFFRX1 \register_reg[5][0]  ( .D(n914), .CK(clk), .RN(n2091), .Q(
        \register[5][0] ) );
  DFFRX1 \register_reg[9][3]  ( .D(n789), .CK(clk), .RN(n2081), .Q(
        \register[9][3] ) );
  DFFRX1 \register_reg[9][2]  ( .D(n788), .CK(clk), .RN(n2081), .Q(
        \register[9][2] ) );
  DFFRX1 \register_reg[9][1]  ( .D(n787), .CK(clk), .RN(n2081), .Q(
        \register[9][1] ) );
  DFFRX1 \register_reg[9][0]  ( .D(n786), .CK(clk), .RN(n2081), .Q(
        \register[9][0] ) );
  DFFRX1 \register_reg[13][3]  ( .D(n661), .CK(clk), .RN(n2071), .Q(
        \register[13][3] ) );
  DFFRX1 \register_reg[13][2]  ( .D(n660), .CK(clk), .RN(n2071), .Q(
        \register[13][2] ) );
  DFFRX1 \register_reg[13][1]  ( .D(n659), .CK(clk), .RN(n2071), .Q(
        \register[13][1] ) );
  DFFRX1 \register_reg[13][0]  ( .D(n658), .CK(clk), .RN(n2071), .Q(
        \register[13][0] ) );
  DFFRX1 \register_reg[17][3]  ( .D(n533), .CK(clk), .RN(n2061), .Q(
        \register[17][3] ) );
  DFFRX1 \register_reg[17][2]  ( .D(n532), .CK(clk), .RN(n2061), .Q(
        \register[17][2] ) );
  DFFRX1 \register_reg[17][1]  ( .D(n531), .CK(clk), .RN(n2061), .Q(
        \register[17][1] ) );
  DFFRX1 \register_reg[17][0]  ( .D(n530), .CK(clk), .RN(n2061), .Q(
        \register[17][0] ) );
  DFFRX1 \register_reg[21][3]  ( .D(n405), .CK(clk), .RN(n2051), .Q(
        \register[21][3] ) );
  DFFRX1 \register_reg[21][2]  ( .D(n404), .CK(clk), .RN(n2051), .Q(
        \register[21][2] ) );
  DFFRX1 \register_reg[21][1]  ( .D(n403), .CK(clk), .RN(n2051), .Q(
        \register[21][1] ) );
  DFFRX1 \register_reg[21][0]  ( .D(n402), .CK(clk), .RN(n2051), .Q(
        \register[21][0] ) );
  DFFRX1 \register_reg[25][2]  ( .D(n276), .CK(clk), .RN(n2041), .Q(
        \register[25][2] ) );
  DFFRX1 \register_reg[25][1]  ( .D(n275), .CK(clk), .RN(n2041), .Q(
        \register[25][1] ) );
  DFFRX1 \register_reg[25][0]  ( .D(n274), .CK(clk), .RN(n2041), .Q(
        \register[25][0] ) );
  DFFRX1 \register_reg[29][2]  ( .D(n148), .CK(clk), .RN(n2032), .Q(
        \register[29][2] ) );
  DFFRX1 \register_reg[29][1]  ( .D(n147), .CK(clk), .RN(n2032), .Q(
        \register[29][1] ) );
  DFFRX1 \register_reg[29][0]  ( .D(n146), .CK(clk), .RN(n2031), .Q(
        \register[29][0] ) );
  DFFRX1 \register_reg[0][3]  ( .D(n1077), .CK(clk), .RN(n2103), .Q(
        \register[0][3] ) );
  DFFRX1 \register_reg[0][2]  ( .D(n1076), .CK(clk), .RN(n2103), .Q(
        \register[0][2] ) );
  DFFRX1 \register_reg[0][1]  ( .D(n1075), .CK(clk), .RN(n2103), .Q(
        \register[0][1] ) );
  DFFRX1 \register_reg[0][0]  ( .D(n1074), .CK(clk), .RN(n2103), .Q(
        \register[0][0] ) );
  DFFRX1 \register_reg[4][3]  ( .D(n949), .CK(clk), .RN(n2093), .Q(
        \register[4][3] ) );
  DFFRX1 \register_reg[4][2]  ( .D(n948), .CK(clk), .RN(n2093), .Q(
        \register[4][2] ) );
  DFFRX1 \register_reg[4][1]  ( .D(n947), .CK(clk), .RN(n2093), .Q(
        \register[4][1] ) );
  DFFRX1 \register_reg[4][0]  ( .D(n946), .CK(clk), .RN(n2093), .Q(
        \register[4][0] ) );
  DFFRX1 \register_reg[8][3]  ( .D(n821), .CK(clk), .RN(n2083), .Q(
        \register[8][3] ) );
  DFFRX1 \register_reg[8][2]  ( .D(n820), .CK(clk), .RN(n2083), .Q(
        \register[8][2] ) );
  DFFRX1 \register_reg[8][1]  ( .D(n819), .CK(clk), .RN(n2083), .Q(
        \register[8][1] ) );
  DFFRX1 \register_reg[8][0]  ( .D(n818), .CK(clk), .RN(n2083), .Q(
        \register[8][0] ) );
  DFFRX1 \register_reg[12][3]  ( .D(n693), .CK(clk), .RN(n2074), .Q(
        \register[12][3] ) );
  DFFRX1 \register_reg[12][2]  ( .D(n692), .CK(clk), .RN(n2073), .Q(
        \register[12][2] ) );
  DFFRX1 \register_reg[12][1]  ( .D(n691), .CK(clk), .RN(n2073), .Q(
        \register[12][1] ) );
  DFFRX1 \register_reg[12][0]  ( .D(n690), .CK(clk), .RN(n2073), .Q(
        \register[12][0] ) );
  DFFRX1 \register_reg[16][3]  ( .D(n565), .CK(clk), .RN(n2064), .Q(
        \register[16][3] ) );
  DFFRX1 \register_reg[16][2]  ( .D(n564), .CK(clk), .RN(n2064), .Q(
        \register[16][2] ) );
  DFFRX1 \register_reg[16][1]  ( .D(n563), .CK(clk), .RN(n2064), .Q(
        \register[16][1] ) );
  DFFRX1 \register_reg[16][0]  ( .D(n562), .CK(clk), .RN(n2063), .Q(
        \register[16][0] ) );
  DFFRX1 \register_reg[20][3]  ( .D(n437), .CK(clk), .RN(n2054), .Q(
        \register[20][3] ) );
  DFFRX1 \register_reg[20][2]  ( .D(n436), .CK(clk), .RN(n2054), .Q(
        \register[20][2] ) );
  DFFRX1 \register_reg[20][1]  ( .D(n435), .CK(clk), .RN(n2054), .Q(
        \register[20][1] ) );
  DFFRX1 \register_reg[20][0]  ( .D(n434), .CK(clk), .RN(n2054), .Q(
        \register[20][0] ) );
  DFFRX1 \register_reg[24][3]  ( .D(n309), .CK(clk), .RN(n2044), .Q(
        \register[24][3] ) );
  DFFRX1 \register_reg[24][2]  ( .D(n308), .CK(clk), .RN(n2044), .Q(
        \register[24][2] ) );
  DFFRX1 \register_reg[24][1]  ( .D(n307), .CK(clk), .RN(n2044), .Q(
        \register[24][1] ) );
  DFFRX1 \register_reg[24][0]  ( .D(n306), .CK(clk), .RN(n2044), .Q(
        \register[24][0] ) );
  DFFRX1 \register_reg[28][2]  ( .D(n180), .CK(clk), .RN(n2034), .Q(
        \register[28][2] ) );
  DFFRX1 \register_reg[28][1]  ( .D(n179), .CK(clk), .RN(n2034), .Q(
        \register[28][1] ) );
  DFFRX1 \register_reg[28][0]  ( .D(n178), .CK(clk), .RN(n2034), .Q(
        \register[28][0] ) );
  DFFRX1 \register_reg[2][3]  ( .D(n1013), .CK(clk), .RN(n2098), .Q(
        \register[2][3] ) );
  DFFRX1 \register_reg[2][2]  ( .D(n1012), .CK(clk), .RN(n2098), .Q(
        \register[2][2] ) );
  DFFRX1 \register_reg[2][1]  ( .D(n1011), .CK(clk), .RN(n2098), .Q(
        \register[2][1] ) );
  DFFRX1 \register_reg[2][0]  ( .D(n1010), .CK(clk), .RN(n2098), .Q(
        \register[2][0] ) );
  DFFRX1 \register_reg[6][3]  ( .D(n885), .CK(clk), .RN(n2088), .Q(
        \register[6][3] ) );
  DFFRX1 \register_reg[6][2]  ( .D(n884), .CK(clk), .RN(n2088), .Q(
        \register[6][2] ) );
  DFFRX1 \register_reg[6][1]  ( .D(n883), .CK(clk), .RN(n2088), .Q(
        \register[6][1] ) );
  DFFRX1 \register_reg[6][0]  ( .D(n882), .CK(clk), .RN(n2088), .Q(
        \register[6][0] ) );
  DFFRX1 \register_reg[10][3]  ( .D(n757), .CK(clk), .RN(n2078), .Q(
        \register[10][3] ) );
  DFFRX1 \register_reg[10][2]  ( .D(n756), .CK(clk), .RN(n2078), .Q(
        \register[10][2] ) );
  DFFRX1 \register_reg[10][1]  ( .D(n755), .CK(clk), .RN(n2078), .Q(
        \register[10][1] ) );
  DFFRX1 \register_reg[10][0]  ( .D(n754), .CK(clk), .RN(n2078), .Q(
        \register[10][0] ) );
  DFFRX1 \register_reg[14][3]  ( .D(n629), .CK(clk), .RN(n2069), .Q(
        \register[14][3] ) );
  DFFRX1 \register_reg[14][2]  ( .D(n628), .CK(clk), .RN(n2069), .Q(
        \register[14][2] ) );
  DFFRX1 \register_reg[14][1]  ( .D(n627), .CK(clk), .RN(n2068), .Q(
        \register[14][1] ) );
  DFFRX1 \register_reg[14][0]  ( .D(n626), .CK(clk), .RN(n2068), .Q(
        \register[14][0] ) );
  DFFRX1 \register_reg[18][3]  ( .D(n501), .CK(clk), .RN(n2059), .Q(
        \register[18][3] ) );
  DFFRX1 \register_reg[18][2]  ( .D(n500), .CK(clk), .RN(n2059), .Q(
        \register[18][2] ) );
  DFFRX1 \register_reg[18][1]  ( .D(n499), .CK(clk), .RN(n2059), .Q(
        \register[18][1] ) );
  DFFRX1 \register_reg[18][0]  ( .D(n498), .CK(clk), .RN(n2059), .Q(
        \register[18][0] ) );
  DFFRX1 \register_reg[22][3]  ( .D(n373), .CK(clk), .RN(n2049), .Q(
        \register[22][3] ) );
  DFFRX1 \register_reg[22][2]  ( .D(n372), .CK(clk), .RN(n2049), .Q(
        \register[22][2] ) );
  DFFRX1 \register_reg[22][1]  ( .D(n371), .CK(clk), .RN(n2049), .Q(
        \register[22][1] ) );
  DFFRX1 \register_reg[22][0]  ( .D(n370), .CK(clk), .RN(n2049), .Q(
        \register[22][0] ) );
  DFFRX1 \register_reg[26][2]  ( .D(n244), .CK(clk), .RN(n2039), .Q(
        \register[26][2] ) );
  DFFRX1 \register_reg[26][1]  ( .D(n243), .CK(clk), .RN(n2039), .Q(
        \register[26][1] ) );
  DFFRX1 \register_reg[26][0]  ( .D(n242), .CK(clk), .RN(n2039), .Q(
        \register[26][0] ) );
  DFFRX1 \register_reg[30][2]  ( .D(n116), .CK(clk), .RN(n2029), .Q(
        \register[30][2] ) );
  DFFRX1 \register_reg[30][1]  ( .D(n115), .CK(clk), .RN(n2029), .Q(
        \register[30][1] ) );
  DFFRX1 \register_reg[30][0]  ( .D(n114), .CK(clk), .RN(n2029), .Q(
        \register[30][0] ) );
  DFFRX1 \register_reg[30][8]  ( .D(n122), .CK(clk), .RN(n2310), .Q(
        \register[30][8] ) );
  DFFRX1 \register_reg[30][7]  ( .D(n121), .CK(clk), .RN(n2310), .Q(
        \register[30][7] ) );
  DFFRX1 \register_reg[30][6]  ( .D(n120), .CK(clk), .RN(n2310), .Q(
        \register[30][6] ) );
  DFFRX1 \register_reg[30][5]  ( .D(n119), .CK(clk), .RN(n2310), .Q(
        \register[30][5] ) );
  DFFRX1 \register_reg[30][4]  ( .D(n118), .CK(clk), .RN(n2310), .Q(
        \register[30][4] ) );
  DFFRX1 \register_reg[30][3]  ( .D(n117), .CK(clk), .RN(n2310), .Q(
        \register[30][3] ) );
  DFFRX1 \register_reg[29][8]  ( .D(n154), .CK(clk), .RN(n2310), .Q(
        \register[29][8] ) );
  DFFRX1 \register_reg[29][7]  ( .D(n153), .CK(clk), .RN(n2310), .Q(
        \register[29][7] ) );
  DFFRX1 \register_reg[29][6]  ( .D(n152), .CK(clk), .RN(n2310), .Q(
        \register[29][6] ) );
  DFFRX1 \register_reg[29][5]  ( .D(n151), .CK(clk), .RN(n2310), .Q(
        \register[29][5] ) );
  DFFRX1 \register_reg[29][4]  ( .D(n150), .CK(clk), .RN(n2310), .Q(
        \register[29][4] ) );
  DFFRX1 \register_reg[29][3]  ( .D(n149), .CK(clk), .RN(n2310), .Q(
        \register[29][3] ) );
  DFFRX1 \register_reg[28][8]  ( .D(n186), .CK(clk), .RN(n2310), .Q(
        \register[28][8] ) );
  DFFRX1 \register_reg[28][7]  ( .D(n185), .CK(clk), .RN(n2310), .Q(
        \register[28][7] ) );
  DFFRX1 \register_reg[28][6]  ( .D(n184), .CK(clk), .RN(n2310), .Q(
        \register[28][6] ) );
  DFFRX1 \register_reg[28][5]  ( .D(n183), .CK(clk), .RN(n2310), .Q(
        \register[28][5] ) );
  DFFRX1 \register_reg[28][4]  ( .D(n182), .CK(clk), .RN(n2310), .Q(
        \register[28][4] ) );
  DFFRX1 \register_reg[28][3]  ( .D(n181), .CK(clk), .RN(n2310), .Q(
        \register[28][3] ) );
  DFFRX1 \register_reg[27][8]  ( .D(n218), .CK(clk), .RN(n2310), .Q(
        \register[27][8] ) );
  DFFRX1 \register_reg[27][7]  ( .D(n217), .CK(clk), .RN(n2310), .Q(
        \register[27][7] ) );
  DFFRX1 \register_reg[27][6]  ( .D(n216), .CK(clk), .RN(n2310), .Q(
        \register[27][6] ) );
  DFFRX1 \register_reg[27][5]  ( .D(n215), .CK(clk), .RN(n2310), .Q(
        \register[27][5] ) );
  DFFRX1 \register_reg[27][4]  ( .D(n214), .CK(clk), .RN(n2310), .Q(
        \register[27][4] ) );
  DFFRX1 \register_reg[27][3]  ( .D(n213), .CK(clk), .RN(n2310), .Q(
        \register[27][3] ) );
  DFFRX1 \register_reg[26][8]  ( .D(n250), .CK(clk), .RN(n2310), .Q(
        \register[26][8] ) );
  DFFRX1 \register_reg[26][7]  ( .D(n249), .CK(clk), .RN(n2310), .Q(
        \register[26][7] ) );
  DFFRX1 \register_reg[26][6]  ( .D(n248), .CK(clk), .RN(n2310), .Q(
        \register[26][6] ) );
  DFFRX1 \register_reg[26][5]  ( .D(n247), .CK(clk), .RN(n2310), .Q(
        \register[26][5] ) );
  DFFRX1 \register_reg[26][4]  ( .D(n246), .CK(clk), .RN(n2310), .Q(
        \register[26][4] ) );
  DFFRX1 \register_reg[26][3]  ( .D(n245), .CK(clk), .RN(n2310), .Q(
        \register[26][3] ) );
  DFFRX1 \register_reg[25][8]  ( .D(n282), .CK(clk), .RN(n2310), .Q(
        \register[25][8] ) );
  DFFRX1 \register_reg[25][7]  ( .D(n281), .CK(clk), .RN(n2310), .Q(
        \register[25][7] ) );
  DFFRX1 \register_reg[25][6]  ( .D(n280), .CK(clk), .RN(n2310), .Q(
        \register[25][6] ) );
  DFFRX1 \register_reg[25][5]  ( .D(n279), .CK(clk), .RN(n2310), .Q(
        \register[25][5] ) );
  DFFRX1 \register_reg[25][4]  ( .D(n278), .CK(clk), .RN(n2310), .Q(
        \register[25][4] ) );
  DFFRX1 \register_reg[25][3]  ( .D(n277), .CK(clk), .RN(n2310), .Q(
        \register[25][3] ) );
  DFFRX1 \register_reg[24][8]  ( .D(n314), .CK(clk), .RN(n2310), .Q(
        \register[24][8] ) );
  DFFRX1 \register_reg[24][7]  ( .D(n313), .CK(clk), .RN(n2310), .Q(
        \register[24][7] ) );
  DFFRX1 \register_reg[24][6]  ( .D(n312), .CK(clk), .RN(n2310), .Q(
        \register[24][6] ) );
  NOR3BXL U2 ( .AN(RegWrite_i), .B(WriteReg_i[4]), .C(n2309), .Y(n65) );
  NOR3BXL U3 ( .AN(RegWrite_i), .B(WriteReg_i[3]), .C(WriteReg_i[4]), .Y(n74)
         );
  INVX3 U4 ( .A(rst), .Y(n2310) );
  NAND2X1 U5 ( .A(n39), .B(n40), .Y(n38) );
  NAND2X1 U6 ( .A(n56), .B(n39), .Y(n55) );
  NAND2X1 U7 ( .A(n65), .B(n39), .Y(n64) );
  NAND2X1 U8 ( .A(n74), .B(n39), .Y(n73) );
  NAND2X1 U9 ( .A(n42), .B(n40), .Y(n41) );
  NAND2X1 U10 ( .A(n44), .B(n40), .Y(n43) );
  NAND2X1 U11 ( .A(n46), .B(n40), .Y(n45) );
  NAND2X1 U12 ( .A(n48), .B(n40), .Y(n47) );
  NAND2X1 U13 ( .A(n50), .B(n40), .Y(n49) );
  NAND2X1 U14 ( .A(n52), .B(n40), .Y(n51) );
  NAND2X1 U15 ( .A(n54), .B(n40), .Y(n53) );
  NAND2X1 U16 ( .A(n56), .B(n54), .Y(n63) );
  NAND2X1 U17 ( .A(n65), .B(n54), .Y(n72) );
  NAND2X1 U18 ( .A(n74), .B(n54), .Y(n81) );
  NAND2X1 U19 ( .A(n65), .B(n42), .Y(n66) );
  NAND2X1 U20 ( .A(n65), .B(n44), .Y(n67) );
  NAND2X1 U21 ( .A(n65), .B(n46), .Y(n68) );
  NAND2X1 U22 ( .A(n65), .B(n48), .Y(n69) );
  NAND2X1 U23 ( .A(n65), .B(n50), .Y(n70) );
  NAND2X1 U24 ( .A(n65), .B(n52), .Y(n71) );
  NAND2X1 U25 ( .A(n56), .B(n42), .Y(n57) );
  NAND2X1 U26 ( .A(n56), .B(n44), .Y(n58) );
  NAND2X1 U27 ( .A(n56), .B(n46), .Y(n59) );
  NAND2X1 U28 ( .A(n74), .B(n42), .Y(n75) );
  NAND2X1 U29 ( .A(n74), .B(n44), .Y(n76) );
  NAND2X1 U30 ( .A(n74), .B(n46), .Y(n77) );
  NAND2X1 U31 ( .A(n56), .B(n48), .Y(n60) );
  NAND2X1 U32 ( .A(n56), .B(n50), .Y(n61) );
  NAND2X1 U33 ( .A(n74), .B(n48), .Y(n78) );
  NAND2X1 U34 ( .A(n74), .B(n50), .Y(n79) );
  NAND2X1 U35 ( .A(n56), .B(n52), .Y(n62) );
  NAND2X1 U36 ( .A(n74), .B(n52), .Y(n80) );
  NOR3X1 U37 ( .A(n2307), .B(WriteReg_i[0]), .C(n2308), .Y(n42) );
  NOR3X1 U38 ( .A(n2306), .B(WriteReg_i[1]), .C(n2308), .Y(n44) );
  NOR3X1 U39 ( .A(WriteReg_i[0]), .B(WriteReg_i[1]), .C(n2308), .Y(n46) );
  NOR3X1 U40 ( .A(n2306), .B(WriteReg_i[2]), .C(n2307), .Y(n48) );
  NOR3X1 U41 ( .A(WriteReg_i[0]), .B(WriteReg_i[2]), .C(n2307), .Y(n50) );
  NOR3X1 U42 ( .A(WriteReg_i[1]), .B(WriteReg_i[2]), .C(n2306), .Y(n52) );
  NOR3X1 U43 ( .A(WriteReg_i[1]), .B(WriteReg_i[2]), .C(WriteReg_i[0]), .Y(n54) );
  CLKINVX1 U44 ( .A(WriteReg_i[2]), .Y(n2308) );
  CLKINVX1 U45 ( .A(WriteReg_i[1]), .Y(n2307) );
  CLKINVX1 U46 ( .A(WriteReg_i[0]), .Y(n2306) );
  MXI2X1 U47 ( .A(n7), .B(n8), .S0(n1389), .Y(ReadData1_o[3]) );
  MXI2X1 U48 ( .A(n3), .B(n4), .S0(n1389), .Y(ReadData1_o[1]) );
  MXI2X1 U49 ( .A(n11), .B(n12), .S0(n1389), .Y(ReadData1_o[5]) );
  MXI2X1 U50 ( .A(n9), .B(n10), .S0(n1389), .Y(ReadData1_o[4]) );
  MXI2X1 U51 ( .A(n5), .B(n6), .S0(n1389), .Y(ReadData1_o[2]) );
  MXI2X1 U52 ( .A(n1), .B(n2), .S0(n1389), .Y(ReadData1_o[0]) );
  MXI2X1 U53 ( .A(n19), .B(n20), .S0(n1390), .Y(ReadData1_o[9]) );
  MXI2X1 U54 ( .A(n17), .B(n18), .S0(n1390), .Y(ReadData1_o[8]) );
  MXI2X1 U55 ( .A(n13), .B(n14), .S0(n1389), .Y(ReadData1_o[6]) );
  MXI2X1 U56 ( .A(n15), .B(n16), .S0(n1389), .Y(ReadData1_o[7]) );
  MXI2X1 U57 ( .A(n23), .B(n24), .S0(n1390), .Y(ReadData1_o[11]) );
  MXI2X1 U58 ( .A(n27), .B(n28), .S0(n1390), .Y(ReadData1_o[13]) );
  MXI2X1 U59 ( .A(n21), .B(n22), .S0(n1390), .Y(ReadData1_o[10]) );
  MXI2X1 U60 ( .A(n25), .B(n26), .S0(n1390), .Y(ReadData1_o[12]) );
  MXI2X1 U61 ( .A(n29), .B(n30), .S0(n1390), .Y(ReadData1_o[14]) );
  MXI2X1 U62 ( .A(n37), .B(n1106), .S0(n1390), .Y(ReadData1_o[18]) );
  MXI2X1 U63 ( .A(n31), .B(n32), .S0(n1390), .Y(ReadData1_o[15]) );
  MXI2X1 U64 ( .A(n33), .B(n34), .S0(n1390), .Y(ReadData1_o[16]) );
  MXI2X1 U65 ( .A(n35), .B(n36), .S0(n1390), .Y(ReadData1_o[17]) );
  MXI2X1 U66 ( .A(n1113), .B(n1114), .S0(n1391), .Y(ReadData1_o[22]) );
  MXI2X1 U67 ( .A(n1111), .B(n1112), .S0(n1391), .Y(ReadData1_o[21]) );
  MXI2X1 U68 ( .A(n1109), .B(n1110), .S0(n1391), .Y(ReadData1_o[20]) );
  MXI2X1 U69 ( .A(n1107), .B(n1108), .S0(n1390), .Y(ReadData1_o[19]) );
  MXI2X1 U70 ( .A(n1121), .B(n1122), .S0(n1391), .Y(ReadData1_o[26]) );
  MXI2X1 U71 ( .A(n1123), .B(n1124), .S0(n1391), .Y(ReadData1_o[27]) );
  MXI2X1 U72 ( .A(n1115), .B(n1116), .S0(n1391), .Y(ReadData1_o[23]) );
  MXI2X1 U73 ( .A(n1119), .B(n1120), .S0(n1391), .Y(ReadData1_o[25]) );
  MXI2X1 U74 ( .A(n1117), .B(n1118), .S0(n1391), .Y(ReadData1_o[24]) );
  MXI2X1 U75 ( .A(n1131), .B(n1132), .S0(n1391), .Y(ReadData1_o[31]) );
  MXI2X1 U76 ( .A(n1127), .B(n1128), .S0(n1391), .Y(ReadData1_o[29]) );
  MXI2X1 U77 ( .A(n1125), .B(n1126), .S0(n1391), .Y(ReadData1_o[28]) );
  MXI2X1 U78 ( .A(n1129), .B(n1130), .S0(n1391), .Y(ReadData1_o[30]) );
  CLKBUFX3 U79 ( .A(n1467), .Y(n1471) );
  CLKBUFX3 U80 ( .A(n1465), .Y(n1475) );
  CLKBUFX3 U81 ( .A(n1465), .Y(n1476) );
  CLKBUFX3 U82 ( .A(n1464), .Y(n1477) );
  CLKBUFX3 U83 ( .A(n1464), .Y(n1478) );
  CLKBUFX3 U84 ( .A(n1463), .Y(n1480) );
  CLKBUFX3 U85 ( .A(n1463), .Y(n1479) );
  CLKBUFX3 U86 ( .A(n1462), .Y(n1481) );
  CLKBUFX3 U87 ( .A(n1462), .Y(n1482) );
  CLKBUFX3 U88 ( .A(n1461), .Y(n1483) );
  CLKBUFX3 U89 ( .A(n1461), .Y(n1484) );
  CLKBUFX3 U90 ( .A(n1460), .Y(n1485) );
  CLKBUFX3 U91 ( .A(n1460), .Y(n1486) );
  CLKBUFX3 U92 ( .A(n1459), .Y(n1487) );
  CLKBUFX3 U93 ( .A(n1459), .Y(n1488) );
  CLKBUFX3 U94 ( .A(n1458), .Y(n1489) );
  CLKBUFX3 U95 ( .A(n1458), .Y(n1490) );
  CLKBUFX3 U96 ( .A(n1467), .Y(n1472) );
  CLKBUFX3 U97 ( .A(n1466), .Y(n1473) );
  CLKBUFX3 U98 ( .A(n1466), .Y(n1474) );
  CLKBUFX3 U99 ( .A(n1891), .Y(n1895) );
  CLKBUFX3 U100 ( .A(n1891), .Y(n1896) );
  CLKBUFX3 U101 ( .A(n1890), .Y(n1897) );
  CLKBUFX3 U102 ( .A(n1890), .Y(n1898) );
  CLKBUFX3 U103 ( .A(n1889), .Y(n1899) );
  CLKBUFX3 U104 ( .A(n1889), .Y(n1900) );
  CLKBUFX3 U105 ( .A(n1888), .Y(n1901) );
  CLKBUFX3 U106 ( .A(n1888), .Y(n1902) );
  CLKBUFX3 U107 ( .A(n1887), .Y(n1903) );
  CLKBUFX3 U108 ( .A(n1887), .Y(n1904) );
  CLKBUFX3 U109 ( .A(n1886), .Y(n1905) );
  CLKBUFX3 U110 ( .A(n1886), .Y(n1906) );
  CLKBUFX3 U111 ( .A(n1885), .Y(n1907) );
  CLKBUFX3 U112 ( .A(n1885), .Y(n1908) );
  CLKBUFX3 U113 ( .A(n1884), .Y(n1909) );
  CLKBUFX3 U114 ( .A(n1884), .Y(n1910) );
  CLKBUFX3 U115 ( .A(n1883), .Y(n1911) );
  CLKBUFX3 U116 ( .A(n1883), .Y(n1912) );
  CLKBUFX3 U117 ( .A(n1882), .Y(n1913) );
  CLKBUFX3 U118 ( .A(n1882), .Y(n1914) );
  CLKBUFX3 U119 ( .A(n1426), .Y(n1430) );
  CLKBUFX3 U120 ( .A(n1424), .Y(n1434) );
  CLKBUFX3 U121 ( .A(n1424), .Y(n1435) );
  CLKBUFX3 U122 ( .A(n1423), .Y(n1436) );
  CLKBUFX3 U123 ( .A(n1423), .Y(n1437) );
  CLKBUFX3 U124 ( .A(n1422), .Y(n1439) );
  CLKBUFX3 U125 ( .A(n1422), .Y(n1438) );
  CLKBUFX3 U126 ( .A(n1421), .Y(n1440) );
  CLKBUFX3 U127 ( .A(n1421), .Y(n1441) );
  CLKBUFX3 U128 ( .A(n1420), .Y(n1442) );
  CLKBUFX3 U129 ( .A(n1420), .Y(n1443) );
  CLKBUFX3 U130 ( .A(n1419), .Y(n1444) );
  CLKBUFX3 U131 ( .A(n1419), .Y(n1445) );
  CLKBUFX3 U132 ( .A(n1418), .Y(n1446) );
  CLKBUFX3 U133 ( .A(n1418), .Y(n1447) );
  CLKBUFX3 U134 ( .A(n1417), .Y(n1448) );
  CLKBUFX3 U135 ( .A(n1417), .Y(n1449) );
  CLKBUFX3 U136 ( .A(n1426), .Y(n1431) );
  CLKBUFX3 U137 ( .A(n1425), .Y(n1432) );
  CLKBUFX3 U138 ( .A(n1425), .Y(n1433) );
  CLKBUFX3 U139 ( .A(n1850), .Y(n1854) );
  CLKBUFX3 U140 ( .A(n1850), .Y(n1855) );
  CLKBUFX3 U141 ( .A(n1849), .Y(n1856) );
  CLKBUFX3 U142 ( .A(n1849), .Y(n1857) );
  CLKBUFX3 U143 ( .A(n1848), .Y(n1858) );
  CLKBUFX3 U144 ( .A(n1848), .Y(n1859) );
  CLKBUFX3 U145 ( .A(n1847), .Y(n1860) );
  CLKBUFX3 U146 ( .A(n1847), .Y(n1861) );
  CLKBUFX3 U147 ( .A(n1846), .Y(n1862) );
  CLKBUFX3 U148 ( .A(n1846), .Y(n1863) );
  CLKBUFX3 U149 ( .A(n1845), .Y(n1864) );
  CLKBUFX3 U150 ( .A(n1845), .Y(n1865) );
  CLKBUFX3 U151 ( .A(n1844), .Y(n1866) );
  CLKBUFX3 U152 ( .A(n1844), .Y(n1867) );
  CLKBUFX3 U153 ( .A(n1843), .Y(n1868) );
  CLKBUFX3 U154 ( .A(n1843), .Y(n1869) );
  CLKBUFX3 U155 ( .A(n1842), .Y(n1870) );
  CLKBUFX3 U156 ( .A(n1842), .Y(n1871) );
  CLKBUFX3 U157 ( .A(n1841), .Y(n1872) );
  CLKBUFX3 U158 ( .A(n1841), .Y(n1873) );
  CLKBUFX3 U159 ( .A(n38), .Y(n2272) );
  CLKBUFX3 U160 ( .A(n2144), .Y(n2028) );
  CLKBUFX3 U161 ( .A(n2144), .Y(n2029) );
  CLKBUFX3 U162 ( .A(n2143), .Y(n2030) );
  CLKBUFX3 U163 ( .A(n2143), .Y(n2031) );
  CLKBUFX3 U164 ( .A(n2142), .Y(n2032) );
  CLKBUFX3 U165 ( .A(n2142), .Y(n2033) );
  CLKBUFX3 U166 ( .A(n2141), .Y(n2034) );
  CLKBUFX3 U167 ( .A(n2141), .Y(n2035) );
  CLKBUFX3 U168 ( .A(n2140), .Y(n2036) );
  CLKBUFX3 U169 ( .A(n2140), .Y(n2037) );
  CLKBUFX3 U170 ( .A(n2139), .Y(n2038) );
  CLKBUFX3 U171 ( .A(n2139), .Y(n2039) );
  CLKBUFX3 U172 ( .A(n2138), .Y(n2040) );
  CLKBUFX3 U173 ( .A(n2138), .Y(n2041) );
  CLKBUFX3 U174 ( .A(n2137), .Y(n2042) );
  CLKBUFX3 U175 ( .A(n2137), .Y(n2043) );
  CLKBUFX3 U176 ( .A(n2136), .Y(n2044) );
  CLKBUFX3 U177 ( .A(n2136), .Y(n2045) );
  CLKBUFX3 U178 ( .A(n2135), .Y(n2046) );
  CLKBUFX3 U179 ( .A(n2135), .Y(n2047) );
  CLKBUFX3 U180 ( .A(n2134), .Y(n2048) );
  CLKBUFX3 U181 ( .A(n2134), .Y(n2049) );
  CLKBUFX3 U182 ( .A(n2133), .Y(n2050) );
  CLKBUFX3 U183 ( .A(n2133), .Y(n2051) );
  CLKBUFX3 U184 ( .A(n2132), .Y(n2052) );
  CLKBUFX3 U185 ( .A(n2132), .Y(n2053) );
  CLKBUFX3 U186 ( .A(n2131), .Y(n2054) );
  CLKBUFX3 U187 ( .A(n2131), .Y(n2055) );
  CLKBUFX3 U188 ( .A(n2130), .Y(n2056) );
  CLKBUFX3 U189 ( .A(n2130), .Y(n2057) );
  CLKBUFX3 U190 ( .A(n2129), .Y(n2058) );
  CLKBUFX3 U191 ( .A(n2129), .Y(n2059) );
  CLKBUFX3 U192 ( .A(n2128), .Y(n2060) );
  CLKBUFX3 U193 ( .A(n2128), .Y(n2061) );
  CLKBUFX3 U194 ( .A(n2127), .Y(n2062) );
  CLKBUFX3 U195 ( .A(n2127), .Y(n2063) );
  CLKBUFX3 U196 ( .A(n2126), .Y(n2064) );
  CLKBUFX3 U197 ( .A(n2126), .Y(n2065) );
  CLKBUFX3 U198 ( .A(n2125), .Y(n2066) );
  CLKBUFX3 U199 ( .A(n2125), .Y(n2067) );
  CLKBUFX3 U200 ( .A(n2124), .Y(n2068) );
  CLKBUFX3 U201 ( .A(n2124), .Y(n2069) );
  CLKBUFX3 U202 ( .A(n2123), .Y(n2070) );
  CLKBUFX3 U203 ( .A(n2123), .Y(n2071) );
  CLKBUFX3 U204 ( .A(n2122), .Y(n2072) );
  CLKBUFX3 U205 ( .A(n2122), .Y(n2073) );
  CLKBUFX3 U206 ( .A(n2121), .Y(n2074) );
  CLKBUFX3 U207 ( .A(n2121), .Y(n2075) );
  CLKBUFX3 U208 ( .A(n2120), .Y(n2076) );
  CLKBUFX3 U209 ( .A(n2120), .Y(n2077) );
  CLKBUFX3 U210 ( .A(n2119), .Y(n2078) );
  CLKBUFX3 U211 ( .A(n2119), .Y(n2079) );
  CLKBUFX3 U212 ( .A(n2118), .Y(n2080) );
  CLKBUFX3 U213 ( .A(n2118), .Y(n2081) );
  CLKBUFX3 U214 ( .A(n2117), .Y(n2082) );
  CLKBUFX3 U215 ( .A(n2117), .Y(n2083) );
  CLKBUFX3 U216 ( .A(n2116), .Y(n2084) );
  CLKBUFX3 U217 ( .A(n2116), .Y(n2085) );
  CLKBUFX3 U218 ( .A(n2115), .Y(n2086) );
  CLKBUFX3 U219 ( .A(n2115), .Y(n2087) );
  CLKBUFX3 U220 ( .A(n2114), .Y(n2088) );
  CLKBUFX3 U221 ( .A(n2114), .Y(n2089) );
  CLKBUFX3 U222 ( .A(n2113), .Y(n2090) );
  CLKBUFX3 U223 ( .A(n2113), .Y(n2091) );
  CLKBUFX3 U224 ( .A(n2112), .Y(n2092) );
  CLKBUFX3 U225 ( .A(n2112), .Y(n2093) );
  CLKBUFX3 U226 ( .A(n2111), .Y(n2094) );
  CLKBUFX3 U227 ( .A(n2111), .Y(n2095) );
  CLKBUFX3 U228 ( .A(n2110), .Y(n2096) );
  CLKBUFX3 U229 ( .A(n2110), .Y(n2097) );
  CLKBUFX3 U230 ( .A(n2109), .Y(n2098) );
  CLKBUFX3 U231 ( .A(n2109), .Y(n2099) );
  CLKBUFX3 U232 ( .A(n2108), .Y(n2100) );
  CLKBUFX3 U233 ( .A(n2108), .Y(n2101) );
  CLKBUFX3 U234 ( .A(n2107), .Y(n2102) );
  CLKBUFX3 U235 ( .A(n2107), .Y(n2103) );
  CLKBUFX3 U236 ( .A(n2106), .Y(n2104) );
  CLKBUFX3 U237 ( .A(n38), .Y(n2271) );
  CLKBUFX3 U238 ( .A(n38), .Y(n2270) );
  CLKBUFX3 U239 ( .A(n64), .Y(n2208) );
  CLKBUFX3 U240 ( .A(n66), .Y(n2204) );
  CLKBUFX3 U241 ( .A(n67), .Y(n2200) );
  CLKBUFX3 U242 ( .A(n68), .Y(n2196) );
  CLKBUFX3 U243 ( .A(n69), .Y(n2192) );
  CLKBUFX3 U244 ( .A(n70), .Y(n2188) );
  CLKBUFX3 U245 ( .A(n71), .Y(n2184) );
  CLKBUFX3 U246 ( .A(n72), .Y(n2180) );
  CLKBUFX3 U247 ( .A(n73), .Y(n2176) );
  CLKBUFX3 U248 ( .A(n75), .Y(n2172) );
  CLKBUFX3 U249 ( .A(n76), .Y(n2168) );
  CLKBUFX3 U250 ( .A(n77), .Y(n2164) );
  CLKBUFX3 U251 ( .A(n78), .Y(n2160) );
  CLKBUFX3 U252 ( .A(n79), .Y(n2156) );
  CLKBUFX3 U253 ( .A(n80), .Y(n2152) );
  CLKBUFX3 U254 ( .A(n81), .Y(n2148) );
  CLKBUFX3 U255 ( .A(n64), .Y(n2207) );
  CLKBUFX3 U256 ( .A(n64), .Y(n2206) );
  CLKBUFX3 U257 ( .A(n66), .Y(n2203) );
  CLKBUFX3 U258 ( .A(n66), .Y(n2202) );
  CLKBUFX3 U259 ( .A(n67), .Y(n2199) );
  CLKBUFX3 U260 ( .A(n67), .Y(n2198) );
  CLKBUFX3 U261 ( .A(n68), .Y(n2195) );
  CLKBUFX3 U262 ( .A(n68), .Y(n2194) );
  CLKBUFX3 U263 ( .A(n69), .Y(n2191) );
  CLKBUFX3 U264 ( .A(n69), .Y(n2190) );
  CLKBUFX3 U265 ( .A(n70), .Y(n2187) );
  CLKBUFX3 U266 ( .A(n70), .Y(n2186) );
  CLKBUFX3 U267 ( .A(n71), .Y(n2183) );
  CLKBUFX3 U268 ( .A(n71), .Y(n2182) );
  CLKBUFX3 U269 ( .A(n72), .Y(n2179) );
  CLKBUFX3 U270 ( .A(n72), .Y(n2178) );
  CLKBUFX3 U271 ( .A(n73), .Y(n2175) );
  CLKBUFX3 U272 ( .A(n73), .Y(n2174) );
  CLKBUFX3 U273 ( .A(n75), .Y(n2171) );
  CLKBUFX3 U274 ( .A(n75), .Y(n2170) );
  CLKBUFX3 U275 ( .A(n76), .Y(n2167) );
  CLKBUFX3 U276 ( .A(n76), .Y(n2166) );
  CLKBUFX3 U277 ( .A(n77), .Y(n2163) );
  CLKBUFX3 U278 ( .A(n77), .Y(n2162) );
  CLKBUFX3 U279 ( .A(n78), .Y(n2159) );
  CLKBUFX3 U280 ( .A(n78), .Y(n2158) );
  CLKBUFX3 U281 ( .A(n79), .Y(n2155) );
  CLKBUFX3 U282 ( .A(n79), .Y(n2154) );
  CLKBUFX3 U283 ( .A(n80), .Y(n2151) );
  CLKBUFX3 U284 ( .A(n80), .Y(n2150) );
  CLKBUFX3 U285 ( .A(n81), .Y(n2147) );
  CLKBUFX3 U286 ( .A(n81), .Y(n2146) );
  CLKBUFX3 U287 ( .A(n41), .Y(n2268) );
  CLKBUFX3 U288 ( .A(n43), .Y(n2264) );
  CLKBUFX3 U289 ( .A(n45), .Y(n2260) );
  CLKBUFX3 U290 ( .A(n47), .Y(n2256) );
  CLKBUFX3 U291 ( .A(n49), .Y(n2252) );
  CLKBUFX3 U292 ( .A(n51), .Y(n2248) );
  CLKBUFX3 U293 ( .A(n53), .Y(n2244) );
  CLKBUFX3 U294 ( .A(n55), .Y(n2240) );
  CLKBUFX3 U295 ( .A(n57), .Y(n2236) );
  CLKBUFX3 U296 ( .A(n58), .Y(n2232) );
  CLKBUFX3 U297 ( .A(n59), .Y(n2228) );
  CLKBUFX3 U298 ( .A(n60), .Y(n2224) );
  CLKBUFX3 U299 ( .A(n61), .Y(n2220) );
  CLKBUFX3 U300 ( .A(n62), .Y(n2216) );
  CLKBUFX3 U301 ( .A(n63), .Y(n2212) );
  CLKBUFX3 U302 ( .A(n41), .Y(n2267) );
  CLKBUFX3 U303 ( .A(n41), .Y(n2266) );
  CLKBUFX3 U304 ( .A(n43), .Y(n2263) );
  CLKBUFX3 U305 ( .A(n43), .Y(n2262) );
  CLKBUFX3 U306 ( .A(n45), .Y(n2259) );
  CLKBUFX3 U307 ( .A(n45), .Y(n2258) );
  CLKBUFX3 U308 ( .A(n47), .Y(n2255) );
  CLKBUFX3 U309 ( .A(n47), .Y(n2254) );
  CLKBUFX3 U310 ( .A(n49), .Y(n2251) );
  CLKBUFX3 U311 ( .A(n49), .Y(n2250) );
  CLKBUFX3 U312 ( .A(n51), .Y(n2247) );
  CLKBUFX3 U313 ( .A(n51), .Y(n2246) );
  CLKBUFX3 U314 ( .A(n53), .Y(n2243) );
  CLKBUFX3 U315 ( .A(n53), .Y(n2242) );
  CLKBUFX3 U316 ( .A(n55), .Y(n2239) );
  CLKBUFX3 U317 ( .A(n55), .Y(n2238) );
  CLKBUFX3 U318 ( .A(n57), .Y(n2235) );
  CLKBUFX3 U319 ( .A(n57), .Y(n2234) );
  CLKBUFX3 U320 ( .A(n58), .Y(n2231) );
  CLKBUFX3 U321 ( .A(n58), .Y(n2230) );
  CLKBUFX3 U322 ( .A(n59), .Y(n2227) );
  CLKBUFX3 U323 ( .A(n59), .Y(n2226) );
  CLKBUFX3 U324 ( .A(n60), .Y(n2223) );
  CLKBUFX3 U325 ( .A(n60), .Y(n2222) );
  CLKBUFX3 U326 ( .A(n61), .Y(n2219) );
  CLKBUFX3 U327 ( .A(n61), .Y(n2218) );
  CLKBUFX3 U328 ( .A(n62), .Y(n2215) );
  CLKBUFX3 U329 ( .A(n62), .Y(n2214) );
  CLKBUFX3 U330 ( .A(n63), .Y(n2211) );
  CLKBUFX3 U331 ( .A(n63), .Y(n2210) );
  CLKBUFX3 U332 ( .A(n2106), .Y(n2105) );
  CLKBUFX3 U333 ( .A(n1468), .Y(n1470) );
  CLKBUFX3 U334 ( .A(n1892), .Y(n1894) );
  CLKBUFX3 U335 ( .A(n64), .Y(n2209) );
  CLKBUFX3 U336 ( .A(n66), .Y(n2205) );
  CLKBUFX3 U337 ( .A(n67), .Y(n2201) );
  CLKBUFX3 U338 ( .A(n68), .Y(n2197) );
  CLKBUFX3 U339 ( .A(n69), .Y(n2193) );
  CLKBUFX3 U340 ( .A(n70), .Y(n2189) );
  CLKBUFX3 U341 ( .A(n71), .Y(n2185) );
  CLKBUFX3 U342 ( .A(n72), .Y(n2181) );
  CLKBUFX3 U343 ( .A(n73), .Y(n2177) );
  CLKBUFX3 U344 ( .A(n75), .Y(n2173) );
  CLKBUFX3 U345 ( .A(n76), .Y(n2169) );
  CLKBUFX3 U346 ( .A(n77), .Y(n2165) );
  CLKBUFX3 U347 ( .A(n78), .Y(n2161) );
  CLKBUFX3 U348 ( .A(n79), .Y(n2157) );
  CLKBUFX3 U349 ( .A(n80), .Y(n2153) );
  CLKBUFX3 U350 ( .A(n81), .Y(n2149) );
  CLKBUFX3 U351 ( .A(n41), .Y(n2269) );
  CLKBUFX3 U352 ( .A(n43), .Y(n2265) );
  CLKBUFX3 U353 ( .A(n45), .Y(n2261) );
  CLKBUFX3 U354 ( .A(n47), .Y(n2257) );
  CLKBUFX3 U355 ( .A(n49), .Y(n2253) );
  CLKBUFX3 U356 ( .A(n51), .Y(n2249) );
  CLKBUFX3 U357 ( .A(n53), .Y(n2245) );
  CLKBUFX3 U358 ( .A(n57), .Y(n2237) );
  CLKBUFX3 U359 ( .A(n58), .Y(n2233) );
  CLKBUFX3 U360 ( .A(n59), .Y(n2229) );
  CLKBUFX3 U361 ( .A(n63), .Y(n2213) );
  CLKBUFX3 U362 ( .A(n60), .Y(n2225) );
  CLKBUFX3 U363 ( .A(n61), .Y(n2221) );
  CLKBUFX3 U364 ( .A(n62), .Y(n2217) );
  CLKBUFX3 U365 ( .A(n55), .Y(n2241) );
  CLKBUFX3 U366 ( .A(n38), .Y(n2273) );
  CLKBUFX3 U367 ( .A(n1453), .Y(n1467) );
  CLKBUFX3 U368 ( .A(n1412), .Y(n1426) );
  CLKBUFX3 U369 ( .A(n1454), .Y(n1465) );
  CLKBUFX3 U370 ( .A(n1413), .Y(n1424) );
  CLKBUFX3 U371 ( .A(n1454), .Y(n1464) );
  CLKBUFX3 U372 ( .A(n1413), .Y(n1423) );
  CLKBUFX3 U373 ( .A(n1455), .Y(n1463) );
  CLKBUFX3 U374 ( .A(n1414), .Y(n1422) );
  CLKBUFX3 U375 ( .A(n1455), .Y(n1462) );
  CLKBUFX3 U376 ( .A(n1414), .Y(n1421) );
  CLKBUFX3 U377 ( .A(n1456), .Y(n1461) );
  CLKBUFX3 U378 ( .A(n1415), .Y(n1420) );
  CLKBUFX3 U379 ( .A(n1456), .Y(n1460) );
  CLKBUFX3 U380 ( .A(n1415), .Y(n1419) );
  CLKBUFX3 U381 ( .A(n1457), .Y(n1459) );
  CLKBUFX3 U382 ( .A(n1416), .Y(n1418) );
  CLKBUFX3 U383 ( .A(n1457), .Y(n1458) );
  CLKBUFX3 U384 ( .A(n1416), .Y(n1417) );
  CLKBUFX3 U385 ( .A(n1453), .Y(n1466) );
  CLKBUFX3 U386 ( .A(n1412), .Y(n1425) );
  CLKBUFX3 U387 ( .A(n1877), .Y(n1891) );
  CLKBUFX3 U388 ( .A(n1836), .Y(n1850) );
  CLKBUFX3 U389 ( .A(n1877), .Y(n1890) );
  CLKBUFX3 U390 ( .A(n1836), .Y(n1849) );
  CLKBUFX3 U391 ( .A(n1878), .Y(n1889) );
  CLKBUFX3 U392 ( .A(n1837), .Y(n1848) );
  CLKBUFX3 U393 ( .A(n1878), .Y(n1888) );
  CLKBUFX3 U394 ( .A(n1837), .Y(n1847) );
  CLKBUFX3 U395 ( .A(n1879), .Y(n1887) );
  CLKBUFX3 U396 ( .A(n1838), .Y(n1846) );
  CLKBUFX3 U397 ( .A(n1879), .Y(n1886) );
  CLKBUFX3 U398 ( .A(n1838), .Y(n1845) );
  CLKBUFX3 U399 ( .A(n1880), .Y(n1885) );
  CLKBUFX3 U400 ( .A(n1839), .Y(n1844) );
  CLKBUFX3 U401 ( .A(n1880), .Y(n1884) );
  CLKBUFX3 U402 ( .A(n1839), .Y(n1843) );
  CLKBUFX3 U403 ( .A(n1881), .Y(n1883) );
  CLKBUFX3 U404 ( .A(n1840), .Y(n1842) );
  CLKBUFX3 U405 ( .A(n1881), .Y(n1882) );
  CLKBUFX3 U406 ( .A(n1840), .Y(n1841) );
  CLKBUFX3 U407 ( .A(n1427), .Y(n1429) );
  CLKBUFX3 U408 ( .A(n1851), .Y(n1853) );
  CLKBUFX3 U409 ( .A(n1468), .Y(n1469) );
  CLKBUFX3 U410 ( .A(n1892), .Y(n1893) );
  CLKBUFX3 U411 ( .A(n1427), .Y(n1428) );
  CLKBUFX3 U412 ( .A(n1851), .Y(n1852) );
  CLKBUFX3 U413 ( .A(n2305), .Y(n2011) );
  CLKBUFX3 U414 ( .A(n2304), .Y(n2008) );
  CLKBUFX3 U415 ( .A(n2303), .Y(n2005) );
  CLKBUFX3 U416 ( .A(n2302), .Y(n2002) );
  CLKBUFX3 U417 ( .A(n2301), .Y(n1999) );
  CLKBUFX3 U418 ( .A(n2300), .Y(n1996) );
  CLKBUFX3 U419 ( .A(n2299), .Y(n1993) );
  CLKBUFX3 U420 ( .A(n2298), .Y(n1990) );
  CLKBUFX3 U421 ( .A(n2297), .Y(n1987) );
  CLKBUFX3 U422 ( .A(n2296), .Y(n1984) );
  CLKBUFX3 U423 ( .A(n2295), .Y(n1981) );
  CLKBUFX3 U424 ( .A(n2294), .Y(n1978) );
  CLKBUFX3 U425 ( .A(n2293), .Y(n1975) );
  CLKBUFX3 U426 ( .A(n2292), .Y(n1972) );
  CLKBUFX3 U427 ( .A(n2291), .Y(n1969) );
  CLKBUFX3 U428 ( .A(n2290), .Y(n1966) );
  CLKBUFX3 U429 ( .A(n2289), .Y(n1963) );
  CLKBUFX3 U430 ( .A(n2288), .Y(n1960) );
  CLKBUFX3 U431 ( .A(n2287), .Y(n1957) );
  CLKBUFX3 U432 ( .A(n2286), .Y(n1954) );
  CLKBUFX3 U433 ( .A(n2285), .Y(n1951) );
  CLKBUFX3 U434 ( .A(n2284), .Y(n1948) );
  CLKBUFX3 U435 ( .A(n2283), .Y(n1945) );
  CLKBUFX3 U436 ( .A(n2282), .Y(n1942) );
  CLKBUFX3 U437 ( .A(n2281), .Y(n1939) );
  CLKBUFX3 U438 ( .A(n2280), .Y(n1936) );
  CLKBUFX3 U439 ( .A(n2279), .Y(n1933) );
  CLKBUFX3 U440 ( .A(n2278), .Y(n1930) );
  CLKBUFX3 U441 ( .A(n2277), .Y(n1927) );
  CLKBUFX3 U442 ( .A(n2276), .Y(n1924) );
  CLKBUFX3 U443 ( .A(n2275), .Y(n1921) );
  CLKBUFX3 U444 ( .A(n2274), .Y(n1918) );
  CLKBUFX3 U445 ( .A(n2305), .Y(n2010) );
  CLKBUFX3 U446 ( .A(n2304), .Y(n2007) );
  CLKBUFX3 U447 ( .A(n2303), .Y(n2004) );
  CLKBUFX3 U448 ( .A(n2302), .Y(n2001) );
  CLKBUFX3 U449 ( .A(n2301), .Y(n1998) );
  CLKBUFX3 U450 ( .A(n2300), .Y(n1995) );
  CLKBUFX3 U451 ( .A(n2299), .Y(n1992) );
  CLKBUFX3 U452 ( .A(n2298), .Y(n1989) );
  CLKBUFX3 U453 ( .A(n2297), .Y(n1986) );
  CLKBUFX3 U454 ( .A(n2296), .Y(n1983) );
  CLKBUFX3 U455 ( .A(n2295), .Y(n1980) );
  CLKBUFX3 U456 ( .A(n2294), .Y(n1977) );
  CLKBUFX3 U457 ( .A(n2293), .Y(n1974) );
  CLKBUFX3 U458 ( .A(n2292), .Y(n1971) );
  CLKBUFX3 U459 ( .A(n2291), .Y(n1968) );
  CLKBUFX3 U460 ( .A(n2290), .Y(n1965) );
  CLKBUFX3 U461 ( .A(n2289), .Y(n1962) );
  CLKBUFX3 U462 ( .A(n2288), .Y(n1959) );
  CLKBUFX3 U463 ( .A(n2287), .Y(n1956) );
  CLKBUFX3 U464 ( .A(n2286), .Y(n1953) );
  CLKBUFX3 U465 ( .A(n2285), .Y(n1950) );
  CLKBUFX3 U466 ( .A(n2284), .Y(n1947) );
  CLKBUFX3 U467 ( .A(n2283), .Y(n1944) );
  CLKBUFX3 U468 ( .A(n2282), .Y(n1941) );
  CLKBUFX3 U469 ( .A(n2281), .Y(n1938) );
  CLKBUFX3 U470 ( .A(n2280), .Y(n1935) );
  CLKBUFX3 U471 ( .A(n2279), .Y(n1932) );
  CLKBUFX3 U472 ( .A(n2278), .Y(n1929) );
  CLKBUFX3 U473 ( .A(n2277), .Y(n1926) );
  CLKBUFX3 U474 ( .A(n2276), .Y(n1923) );
  CLKBUFX3 U475 ( .A(n2275), .Y(n1920) );
  CLKBUFX3 U476 ( .A(n2274), .Y(n1917) );
  CLKBUFX3 U477 ( .A(n2305), .Y(n2012) );
  CLKBUFX3 U478 ( .A(n2304), .Y(n2009) );
  CLKBUFX3 U479 ( .A(n2303), .Y(n2006) );
  CLKBUFX3 U480 ( .A(n2302), .Y(n2003) );
  CLKBUFX3 U481 ( .A(n2301), .Y(n2000) );
  CLKBUFX3 U482 ( .A(n2300), .Y(n1997) );
  CLKBUFX3 U483 ( .A(n2299), .Y(n1994) );
  CLKBUFX3 U484 ( .A(n2298), .Y(n1991) );
  CLKBUFX3 U485 ( .A(n2297), .Y(n1988) );
  CLKBUFX3 U486 ( .A(n2296), .Y(n1985) );
  CLKBUFX3 U487 ( .A(n2295), .Y(n1982) );
  CLKBUFX3 U488 ( .A(n2294), .Y(n1979) );
  CLKBUFX3 U489 ( .A(n2293), .Y(n1976) );
  CLKBUFX3 U490 ( .A(n2292), .Y(n1973) );
  CLKBUFX3 U491 ( .A(n2291), .Y(n1970) );
  CLKBUFX3 U492 ( .A(n2290), .Y(n1967) );
  CLKBUFX3 U493 ( .A(n2289), .Y(n1964) );
  CLKBUFX3 U494 ( .A(n2288), .Y(n1961) );
  CLKBUFX3 U495 ( .A(n2287), .Y(n1958) );
  CLKBUFX3 U496 ( .A(n2286), .Y(n1955) );
  CLKBUFX3 U497 ( .A(n2285), .Y(n1952) );
  CLKBUFX3 U498 ( .A(n2284), .Y(n1949) );
  CLKBUFX3 U499 ( .A(n2283), .Y(n1946) );
  CLKBUFX3 U500 ( .A(n2282), .Y(n1943) );
  CLKBUFX3 U501 ( .A(n2281), .Y(n1940) );
  CLKBUFX3 U502 ( .A(n2280), .Y(n1937) );
  CLKBUFX3 U503 ( .A(n2279), .Y(n1934) );
  CLKBUFX3 U504 ( .A(n2278), .Y(n1931) );
  CLKBUFX3 U505 ( .A(n2277), .Y(n1928) );
  CLKBUFX3 U506 ( .A(n2276), .Y(n1925) );
  CLKBUFX3 U507 ( .A(n2275), .Y(n1922) );
  CLKBUFX3 U508 ( .A(n2274), .Y(n1919) );
  NOR3X1 U509 ( .A(n2307), .B(n2306), .C(n2308), .Y(n39) );
  CLKBUFX3 U510 ( .A(n1401), .Y(n1396) );
  CLKBUFX3 U511 ( .A(n1401), .Y(n1397) );
  CLKBUFX3 U512 ( .A(n1402), .Y(n1398) );
  CLKBUFX3 U513 ( .A(n1402), .Y(n1399) );
  CLKBUFX3 U514 ( .A(n1400), .Y(n1395) );
  CLKBUFX3 U515 ( .A(n1824), .Y(n1819) );
  CLKBUFX3 U516 ( .A(n1825), .Y(n1820) );
  CLKBUFX3 U517 ( .A(n1825), .Y(n1821) );
  CLKBUFX3 U518 ( .A(n1826), .Y(n1822) );
  CLKBUFX3 U519 ( .A(n1826), .Y(n1823) );
  CLKBUFX3 U520 ( .A(n1833), .Y(n1828) );
  CLKBUFX3 U521 ( .A(n1833), .Y(n1829) );
  CLKBUFX3 U522 ( .A(n1834), .Y(n1830) );
  CLKBUFX3 U523 ( .A(n1834), .Y(n1831) );
  CLKBUFX3 U524 ( .A(n1400), .Y(n1394) );
  CLKBUFX3 U525 ( .A(n1824), .Y(n1818) );
  CLKBUFX3 U526 ( .A(n1491), .Y(n1453) );
  CLKBUFX3 U527 ( .A(n1450), .Y(n1412) );
  CLKBUFX3 U528 ( .A(n1491), .Y(n1454) );
  CLKBUFX3 U529 ( .A(n1450), .Y(n1413) );
  CLKBUFX3 U530 ( .A(n1492), .Y(n1455) );
  CLKBUFX3 U531 ( .A(n1451), .Y(n1414) );
  CLKBUFX3 U532 ( .A(n1492), .Y(n1456) );
  CLKBUFX3 U533 ( .A(n1451), .Y(n1415) );
  CLKBUFX3 U534 ( .A(n1492), .Y(n1457) );
  CLKBUFX3 U535 ( .A(n1451), .Y(n1416) );
  CLKBUFX3 U536 ( .A(n1915), .Y(n1877) );
  CLKBUFX3 U537 ( .A(n1874), .Y(n1836) );
  CLKBUFX3 U538 ( .A(n1915), .Y(n1878) );
  CLKBUFX3 U539 ( .A(n1874), .Y(n1837) );
  CLKBUFX3 U540 ( .A(n1916), .Y(n1879) );
  CLKBUFX3 U541 ( .A(n1875), .Y(n1838) );
  CLKBUFX3 U542 ( .A(n1916), .Y(n1880) );
  CLKBUFX3 U543 ( .A(n1875), .Y(n1839) );
  CLKBUFX3 U544 ( .A(n1916), .Y(n1881) );
  CLKBUFX3 U545 ( .A(n1875), .Y(n1840) );
  CLKBUFX3 U546 ( .A(n2025), .Y(n2144) );
  CLKBUFX3 U547 ( .A(n2025), .Y(n2143) );
  CLKBUFX3 U548 ( .A(n2025), .Y(n2142) );
  CLKBUFX3 U549 ( .A(n2024), .Y(n2141) );
  CLKBUFX3 U550 ( .A(n2024), .Y(n2140) );
  CLKBUFX3 U551 ( .A(n2024), .Y(n2139) );
  CLKBUFX3 U552 ( .A(n2023), .Y(n2138) );
  CLKBUFX3 U553 ( .A(n2023), .Y(n2137) );
  CLKBUFX3 U554 ( .A(n2023), .Y(n2136) );
  CLKBUFX3 U555 ( .A(n2022), .Y(n2135) );
  CLKBUFX3 U556 ( .A(n2022), .Y(n2134) );
  CLKBUFX3 U557 ( .A(n2022), .Y(n2133) );
  CLKBUFX3 U558 ( .A(n2021), .Y(n2132) );
  CLKBUFX3 U559 ( .A(n2021), .Y(n2131) );
  CLKBUFX3 U560 ( .A(n2021), .Y(n2130) );
  CLKBUFX3 U561 ( .A(n2020), .Y(n2129) );
  CLKBUFX3 U562 ( .A(n2020), .Y(n2128) );
  CLKBUFX3 U563 ( .A(n2020), .Y(n2127) );
  CLKBUFX3 U564 ( .A(n2019), .Y(n2126) );
  CLKBUFX3 U565 ( .A(n2019), .Y(n2125) );
  CLKBUFX3 U566 ( .A(n2019), .Y(n2124) );
  CLKBUFX3 U567 ( .A(n2018), .Y(n2123) );
  CLKBUFX3 U568 ( .A(n2018), .Y(n2122) );
  CLKBUFX3 U569 ( .A(n2018), .Y(n2121) );
  CLKBUFX3 U570 ( .A(n2017), .Y(n2120) );
  CLKBUFX3 U571 ( .A(n2017), .Y(n2119) );
  CLKBUFX3 U572 ( .A(n2017), .Y(n2118) );
  CLKBUFX3 U573 ( .A(n2016), .Y(n2117) );
  CLKBUFX3 U574 ( .A(n2016), .Y(n2116) );
  CLKBUFX3 U575 ( .A(n2016), .Y(n2115) );
  CLKBUFX3 U576 ( .A(n2015), .Y(n2114) );
  CLKBUFX3 U577 ( .A(n2015), .Y(n2113) );
  CLKBUFX3 U578 ( .A(n2015), .Y(n2112) );
  CLKBUFX3 U579 ( .A(n2014), .Y(n2111) );
  CLKBUFX3 U580 ( .A(n2014), .Y(n2110) );
  CLKBUFX3 U581 ( .A(n2014), .Y(n2109) );
  CLKBUFX3 U582 ( .A(n2013), .Y(n2108) );
  CLKBUFX3 U583 ( .A(n2013), .Y(n2107) );
  CLKBUFX3 U584 ( .A(n2013), .Y(n2106) );
  CLKBUFX3 U585 ( .A(n1452), .Y(n1468) );
  CLKBUFX3 U586 ( .A(n1491), .Y(n1452) );
  CLKBUFX3 U587 ( .A(n1411), .Y(n1427) );
  CLKBUFX3 U588 ( .A(n1450), .Y(n1411) );
  CLKBUFX3 U589 ( .A(n1876), .Y(n1892) );
  CLKBUFX3 U590 ( .A(n1915), .Y(n1876) );
  CLKBUFX3 U591 ( .A(n1835), .Y(n1851) );
  CLKBUFX3 U592 ( .A(n1874), .Y(n1835) );
  CLKINVX1 U593 ( .A(WriteData_i[0]), .Y(n2305) );
  CLKINVX1 U594 ( .A(WriteData_i[1]), .Y(n2304) );
  CLKINVX1 U595 ( .A(WriteData_i[2]), .Y(n2303) );
  CLKINVX1 U596 ( .A(WriteData_i[3]), .Y(n2302) );
  CLKINVX1 U597 ( .A(WriteData_i[4]), .Y(n2301) );
  CLKINVX1 U598 ( .A(WriteData_i[5]), .Y(n2300) );
  CLKINVX1 U599 ( .A(WriteData_i[6]), .Y(n2299) );
  CLKINVX1 U600 ( .A(WriteData_i[7]), .Y(n2298) );
  CLKINVX1 U601 ( .A(WriteData_i[8]), .Y(n2297) );
  CLKINVX1 U602 ( .A(WriteData_i[9]), .Y(n2296) );
  CLKINVX1 U603 ( .A(WriteData_i[10]), .Y(n2295) );
  CLKINVX1 U604 ( .A(WriteData_i[11]), .Y(n2294) );
  CLKINVX1 U605 ( .A(WriteData_i[12]), .Y(n2293) );
  CLKINVX1 U606 ( .A(WriteData_i[13]), .Y(n2292) );
  CLKINVX1 U607 ( .A(WriteData_i[14]), .Y(n2291) );
  CLKINVX1 U608 ( .A(WriteData_i[15]), .Y(n2290) );
  CLKINVX1 U609 ( .A(WriteData_i[16]), .Y(n2289) );
  CLKINVX1 U610 ( .A(WriteData_i[17]), .Y(n2288) );
  CLKINVX1 U611 ( .A(WriteData_i[18]), .Y(n2287) );
  CLKINVX1 U612 ( .A(WriteData_i[19]), .Y(n2286) );
  CLKINVX1 U613 ( .A(WriteData_i[20]), .Y(n2285) );
  CLKINVX1 U614 ( .A(WriteData_i[21]), .Y(n2284) );
  CLKINVX1 U615 ( .A(WriteData_i[22]), .Y(n2283) );
  CLKINVX1 U616 ( .A(WriteData_i[23]), .Y(n2282) );
  CLKINVX1 U617 ( .A(WriteData_i[24]), .Y(n2281) );
  CLKINVX1 U618 ( .A(WriteData_i[25]), .Y(n2280) );
  CLKINVX1 U619 ( .A(WriteData_i[26]), .Y(n2279) );
  CLKINVX1 U620 ( .A(WriteData_i[27]), .Y(n2278) );
  CLKINVX1 U621 ( .A(WriteData_i[28]), .Y(n2277) );
  CLKINVX1 U622 ( .A(WriteData_i[29]), .Y(n2276) );
  CLKINVX1 U623 ( .A(WriteData_i[30]), .Y(n2275) );
  CLKINVX1 U624 ( .A(WriteData_i[31]), .Y(n2274) );
  AND3X2 U625 ( .A(RegWrite_i), .B(n2309), .C(WriteReg_i[4]), .Y(n56) );
  AND3X2 U626 ( .A(RegWrite_i), .B(WriteReg_i[3]), .C(WriteReg_i[4]), .Y(n40)
         );
  CLKBUFX3 U627 ( .A(n1393), .Y(n1390) );
  CLKBUFX3 U628 ( .A(n1393), .Y(n1391) );
  CLKBUFX3 U629 ( .A(n1817), .Y(n1814) );
  CLKBUFX3 U630 ( .A(n1817), .Y(n1815) );
  CLKBUFX3 U631 ( .A(n2145), .Y(n2027) );
  CLKBUFX3 U632 ( .A(n2026), .Y(n2145) );
  CLKBUFX3 U633 ( .A(n2310), .Y(n2026) );
  CLKINVX1 U634 ( .A(WriteReg_i[3]), .Y(n2309) );
  CLKBUFX3 U635 ( .A(n1409), .Y(n1405) );
  CLKBUFX3 U636 ( .A(n1410), .Y(n1406) );
  CLKBUFX3 U637 ( .A(n1410), .Y(n1407) );
  CLKBUFX3 U638 ( .A(n1409), .Y(n1404) );
  CLKBUFX3 U639 ( .A(n1832), .Y(n1827) );
  CLKBUFX3 U640 ( .A(N17), .Y(n1832) );
  CLKBUFX3 U641 ( .A(N13), .Y(n1401) );
  CLKBUFX3 U642 ( .A(N13), .Y(n1402) );
  CLKBUFX3 U643 ( .A(N13), .Y(n1400) );
  CLKBUFX3 U644 ( .A(N18), .Y(n1824) );
  CLKBUFX3 U645 ( .A(N17), .Y(n1833) );
  CLKBUFX3 U646 ( .A(N18), .Y(n1825) );
  CLKBUFX3 U647 ( .A(N18), .Y(n1826) );
  CLKBUFX3 U648 ( .A(N17), .Y(n1834) );
  CLKBUFX3 U649 ( .A(N10), .Y(n1491) );
  CLKBUFX3 U650 ( .A(N11), .Y(n1450) );
  CLKBUFX3 U651 ( .A(N10), .Y(n1492) );
  CLKBUFX3 U652 ( .A(N11), .Y(n1451) );
  CLKBUFX3 U653 ( .A(N15), .Y(n1915) );
  CLKBUFX3 U654 ( .A(N16), .Y(n1874) );
  CLKBUFX3 U655 ( .A(N15), .Y(n1916) );
  CLKBUFX3 U656 ( .A(N16), .Y(n1875) );
  CLKBUFX3 U657 ( .A(n2310), .Y(n2025) );
  CLKBUFX3 U658 ( .A(n2310), .Y(n2024) );
  CLKBUFX3 U659 ( .A(n2310), .Y(n2023) );
  CLKBUFX3 U660 ( .A(n2310), .Y(n2022) );
  CLKBUFX3 U661 ( .A(n2310), .Y(n2021) );
  CLKBUFX3 U662 ( .A(n2310), .Y(n2020) );
  CLKBUFX3 U663 ( .A(n2310), .Y(n2019) );
  CLKBUFX3 U664 ( .A(n2310), .Y(n2018) );
  CLKBUFX3 U665 ( .A(n2310), .Y(n2017) );
  CLKBUFX3 U666 ( .A(n2310), .Y(n2016) );
  CLKBUFX3 U667 ( .A(n2310), .Y(n2015) );
  CLKBUFX3 U668 ( .A(n2310), .Y(n2014) );
  CLKBUFX3 U669 ( .A(n2310), .Y(n2013) );
  MXI2X1 U670 ( .A(n1493), .B(n1494), .S0(n1813), .Y(ReadData2_o[0]) );
  MX4X1 U671 ( .A(n1564), .B(n1562), .C(n1563), .D(n1561), .S0(n1818), .S1(
        n1827), .Y(n1493) );
  MX4X1 U672 ( .A(n1560), .B(n1558), .C(n1559), .D(n1557), .S0(n1818), .S1(
        n1827), .Y(n1494) );
  MXI4X1 U673 ( .A(\register[0][0] ), .B(\register[1][0] ), .C(
        \register[2][0] ), .D(\register[3][0] ), .S0(n1894), .S1(n1853), .Y(
        n1564) );
  MXI2X1 U674 ( .A(n1495), .B(n1496), .S0(n1813), .Y(ReadData2_o[1]) );
  MX4X1 U675 ( .A(n1572), .B(n1570), .C(n1571), .D(n1569), .S0(n1818), .S1(
        n1827), .Y(n1495) );
  MX4X1 U676 ( .A(n1568), .B(n1566), .C(n1567), .D(n1565), .S0(n1818), .S1(
        n1827), .Y(n1496) );
  MXI4X1 U677 ( .A(\register[0][1] ), .B(\register[1][1] ), .C(
        \register[2][1] ), .D(\register[3][1] ), .S0(n1894), .S1(n1853), .Y(
        n1572) );
  MXI2X1 U678 ( .A(n1497), .B(n1498), .S0(n1813), .Y(ReadData2_o[2]) );
  MX4X1 U679 ( .A(n1580), .B(n1578), .C(n1579), .D(n1577), .S0(n1819), .S1(
        n1827), .Y(n1497) );
  MX4X1 U680 ( .A(n1576), .B(n1574), .C(n1575), .D(n1573), .S0(n1819), .S1(
        n1827), .Y(n1498) );
  MXI4X1 U681 ( .A(\register[0][2] ), .B(\register[1][2] ), .C(
        \register[2][2] ), .D(\register[3][2] ), .S0(n1895), .S1(n1854), .Y(
        n1580) );
  MXI2X1 U682 ( .A(n1499), .B(n1500), .S0(n1813), .Y(ReadData2_o[3]) );
  MX4X1 U683 ( .A(n1588), .B(n1586), .C(n1587), .D(n1585), .S0(n1819), .S1(
        n1827), .Y(n1499) );
  MX4X1 U684 ( .A(n1584), .B(n1582), .C(n1583), .D(n1581), .S0(n1819), .S1(
        n1827), .Y(n1500) );
  MXI4X1 U685 ( .A(\register[0][3] ), .B(\register[1][3] ), .C(
        \register[2][3] ), .D(\register[3][3] ), .S0(n1896), .S1(n1855), .Y(
        n1588) );
  MX4X1 U686 ( .A(n1152), .B(n1150), .C(n1151), .D(n1149), .S0(n1395), .S1(
        n1403), .Y(n6) );
  MX4X1 U687 ( .A(n1156), .B(n1154), .C(n1155), .D(n1153), .S0(n1395), .S1(
        n1403), .Y(n5) );
  MXI4X1 U688 ( .A(\register[28][2] ), .B(\register[29][2] ), .C(
        \register[30][2] ), .D(\register[31][2] ), .S0(n1471), .S1(n1430), .Y(
        n1149) );
  MX4X1 U689 ( .A(n1160), .B(n1158), .C(n1159), .D(n1157), .S0(n1395), .S1(
        n1403), .Y(n8) );
  MX4X1 U690 ( .A(n1164), .B(n1162), .C(n1163), .D(n1161), .S0(n1395), .S1(
        n1403), .Y(n7) );
  MXI4X1 U691 ( .A(\register[28][3] ), .B(\register[29][3] ), .C(
        \register[30][3] ), .D(\register[31][3] ), .S0(n1471), .S1(n1430), .Y(
        n1157) );
  MX4X1 U692 ( .A(n1144), .B(n1142), .C(n1143), .D(n1141), .S0(n1394), .S1(
        n1403), .Y(n4) );
  MX4X1 U693 ( .A(n1148), .B(n1146), .C(n1147), .D(n1145), .S0(n1394), .S1(
        n1403), .Y(n3) );
  MXI4X1 U694 ( .A(\register[28][1] ), .B(\register[29][1] ), .C(
        \register[30][1] ), .D(\register[31][1] ), .S0(n1470), .S1(n1429), .Y(
        n1141) );
  MX4X1 U695 ( .A(n1136), .B(n1134), .C(n1135), .D(n1133), .S0(n1394), .S1(
        n1403), .Y(n2) );
  MX4X1 U696 ( .A(n1140), .B(n1138), .C(n1139), .D(n1137), .S0(n1394), .S1(
        n1403), .Y(n1) );
  MXI4X1 U697 ( .A(\register[28][0] ), .B(\register[29][0] ), .C(
        \register[30][0] ), .D(\register[31][0] ), .S0(n1469), .S1(n1428), .Y(
        n1133) );
  MXI4X1 U698 ( .A(\register[20][0] ), .B(\register[21][0] ), .C(
        \register[22][0] ), .D(\register[23][0] ), .S0(n1469), .S1(n1428), .Y(
        n1135) );
  MXI4X1 U699 ( .A(\register[20][0] ), .B(\register[21][0] ), .C(
        \register[22][0] ), .D(\register[23][0] ), .S0(n1893), .S1(n1852), .Y(
        n1559) );
  MXI4X1 U700 ( .A(\register[4][2] ), .B(\register[5][2] ), .C(
        \register[6][2] ), .D(\register[7][2] ), .S0(n1471), .S1(n1430), .Y(
        n1155) );
  MXI4X1 U701 ( .A(\register[20][2] ), .B(\register[21][2] ), .C(
        \register[22][2] ), .D(\register[23][2] ), .S0(n1471), .S1(n1430), .Y(
        n1151) );
  MXI4X1 U702 ( .A(\register[4][3] ), .B(\register[5][3] ), .C(
        \register[6][3] ), .D(\register[7][3] ), .S0(n1472), .S1(n1431), .Y(
        n1163) );
  MXI4X1 U703 ( .A(\register[20][3] ), .B(\register[21][3] ), .C(
        \register[22][3] ), .D(\register[23][3] ), .S0(n1471), .S1(n1430), .Y(
        n1159) );
  MXI4X1 U704 ( .A(\register[4][1] ), .B(\register[5][1] ), .C(
        \register[6][1] ), .D(\register[7][1] ), .S0(n1470), .S1(n1429), .Y(
        n1147) );
  MXI4X1 U705 ( .A(\register[20][1] ), .B(\register[21][1] ), .C(
        \register[22][1] ), .D(\register[23][1] ), .S0(n1470), .S1(n1429), .Y(
        n1143) );
  MXI4X1 U706 ( .A(\register[4][0] ), .B(\register[5][0] ), .C(
        \register[6][0] ), .D(\register[7][0] ), .S0(n1470), .S1(n1429), .Y(
        n1139) );
  MXI4X1 U707 ( .A(\register[4][0] ), .B(\register[5][0] ), .C(
        \register[6][0] ), .D(\register[7][0] ), .S0(n1894), .S1(n1853), .Y(
        n1563) );
  MXI4X1 U708 ( .A(\register[20][1] ), .B(\register[21][1] ), .C(
        \register[22][1] ), .D(\register[23][1] ), .S0(n1894), .S1(n1853), .Y(
        n1567) );
  MXI4X1 U709 ( .A(\register[4][1] ), .B(\register[5][1] ), .C(
        \register[6][1] ), .D(\register[7][1] ), .S0(n1894), .S1(n1853), .Y(
        n1571) );
  MXI4X1 U710 ( .A(\register[20][2] ), .B(\register[21][2] ), .C(
        \register[22][2] ), .D(\register[23][2] ), .S0(n1895), .S1(n1854), .Y(
        n1575) );
  MXI4X1 U711 ( .A(\register[4][2] ), .B(\register[5][2] ), .C(
        \register[6][2] ), .D(\register[7][2] ), .S0(n1895), .S1(n1854), .Y(
        n1579) );
  MXI4X1 U712 ( .A(\register[20][3] ), .B(\register[21][3] ), .C(
        \register[22][3] ), .D(\register[23][3] ), .S0(n1895), .S1(n1854), .Y(
        n1583) );
  MXI4X1 U713 ( .A(\register[4][3] ), .B(\register[5][3] ), .C(
        \register[6][3] ), .D(\register[7][3] ), .S0(n1896), .S1(n1855), .Y(
        n1587) );
  MXI4X1 U714 ( .A(\register[16][0] ), .B(\register[17][0] ), .C(
        \register[18][0] ), .D(\register[19][0] ), .S0(n1469), .S1(n1428), .Y(
        n1136) );
  MXI4X1 U715 ( .A(\register[16][0] ), .B(\register[17][0] ), .C(
        \register[18][0] ), .D(\register[19][0] ), .S0(n1893), .S1(n1852), .Y(
        n1560) );
  MXI4X1 U716 ( .A(\register[0][2] ), .B(\register[1][2] ), .C(
        \register[2][2] ), .D(\register[3][2] ), .S0(n1471), .S1(n1430), .Y(
        n1156) );
  MXI4X1 U717 ( .A(\register[16][2] ), .B(\register[17][2] ), .C(
        \register[18][2] ), .D(\register[19][2] ), .S0(n1471), .S1(n1430), .Y(
        n1152) );
  MXI4X1 U718 ( .A(\register[0][3] ), .B(\register[1][3] ), .C(
        \register[2][3] ), .D(\register[3][3] ), .S0(n1472), .S1(n1431), .Y(
        n1164) );
  MXI4X1 U719 ( .A(\register[16][3] ), .B(\register[17][3] ), .C(
        \register[18][3] ), .D(\register[19][3] ), .S0(n1471), .S1(n1430), .Y(
        n1160) );
  MXI4X1 U720 ( .A(\register[0][1] ), .B(\register[1][1] ), .C(
        \register[2][1] ), .D(\register[3][1] ), .S0(n1470), .S1(n1429), .Y(
        n1148) );
  MXI4X1 U721 ( .A(\register[16][1] ), .B(\register[17][1] ), .C(
        \register[18][1] ), .D(\register[19][1] ), .S0(n1470), .S1(n1429), .Y(
        n1144) );
  MXI4X1 U722 ( .A(\register[0][0] ), .B(\register[1][0] ), .C(
        \register[2][0] ), .D(\register[3][0] ), .S0(n1470), .S1(n1429), .Y(
        n1140) );
  MXI4X1 U723 ( .A(\register[16][1] ), .B(\register[17][1] ), .C(
        \register[18][1] ), .D(\register[19][1] ), .S0(n1894), .S1(n1853), .Y(
        n1568) );
  MXI4X1 U724 ( .A(\register[16][2] ), .B(\register[17][2] ), .C(
        \register[18][2] ), .D(\register[19][2] ), .S0(n1895), .S1(n1854), .Y(
        n1576) );
  MXI4X1 U725 ( .A(\register[16][3] ), .B(\register[17][3] ), .C(
        \register[18][3] ), .D(\register[19][3] ), .S0(n1895), .S1(n1854), .Y(
        n1584) );
  MXI4X1 U726 ( .A(\register[28][0] ), .B(\register[29][0] ), .C(
        \register[30][0] ), .D(\register[31][0] ), .S0(n1893), .S1(n1852), .Y(
        n1557) );
  MXI4X1 U727 ( .A(\register[12][2] ), .B(\register[13][2] ), .C(
        \register[14][2] ), .D(\register[15][2] ), .S0(n1471), .S1(n1430), .Y(
        n1153) );
  MXI4X1 U728 ( .A(\register[12][3] ), .B(\register[13][3] ), .C(
        \register[14][3] ), .D(\register[15][3] ), .S0(n1472), .S1(n1431), .Y(
        n1161) );
  MXI4X1 U729 ( .A(\register[12][1] ), .B(\register[13][1] ), .C(
        \register[14][1] ), .D(\register[15][1] ), .S0(n1470), .S1(n1429), .Y(
        n1145) );
  MXI4X1 U730 ( .A(\register[12][0] ), .B(\register[13][0] ), .C(
        \register[14][0] ), .D(\register[15][0] ), .S0(n1470), .S1(n1429), .Y(
        n1137) );
  MXI4X1 U731 ( .A(\register[12][0] ), .B(\register[13][0] ), .C(
        \register[14][0] ), .D(\register[15][0] ), .S0(n1894), .S1(n1853), .Y(
        n1561) );
  MXI4X1 U732 ( .A(\register[28][1] ), .B(\register[29][1] ), .C(
        \register[30][1] ), .D(\register[31][1] ), .S0(n1894), .S1(n1853), .Y(
        n1565) );
  MXI4X1 U733 ( .A(\register[12][1] ), .B(\register[13][1] ), .C(
        \register[14][1] ), .D(\register[15][1] ), .S0(n1894), .S1(n1853), .Y(
        n1569) );
  MXI4X1 U734 ( .A(\register[28][2] ), .B(\register[29][2] ), .C(
        \register[30][2] ), .D(\register[31][2] ), .S0(n1895), .S1(n1854), .Y(
        n1573) );
  MXI4X1 U735 ( .A(\register[12][2] ), .B(\register[13][2] ), .C(
        \register[14][2] ), .D(\register[15][2] ), .S0(n1895), .S1(n1854), .Y(
        n1577) );
  MXI4X1 U736 ( .A(\register[28][3] ), .B(\register[29][3] ), .C(
        \register[30][3] ), .D(\register[31][3] ), .S0(n1895), .S1(n1854), .Y(
        n1581) );
  MXI4X1 U737 ( .A(\register[12][3] ), .B(\register[13][3] ), .C(
        \register[14][3] ), .D(\register[15][3] ), .S0(n1896), .S1(n1855), .Y(
        n1585) );
  MXI4X1 U738 ( .A(\register[24][0] ), .B(\register[25][0] ), .C(
        \register[26][0] ), .D(\register[27][0] ), .S0(n1469), .S1(n1428), .Y(
        n1134) );
  MXI4X1 U739 ( .A(\register[24][0] ), .B(\register[25][0] ), .C(
        \register[26][0] ), .D(\register[27][0] ), .S0(n1893), .S1(n1852), .Y(
        n1558) );
  MXI4X1 U740 ( .A(\register[8][2] ), .B(\register[9][2] ), .C(
        \register[10][2] ), .D(\register[11][2] ), .S0(n1471), .S1(n1430), .Y(
        n1154) );
  MXI4X1 U741 ( .A(\register[24][2] ), .B(\register[25][2] ), .C(
        \register[26][2] ), .D(\register[27][2] ), .S0(n1471), .S1(n1430), .Y(
        n1150) );
  MXI4X1 U742 ( .A(\register[8][3] ), .B(\register[9][3] ), .C(
        \register[10][3] ), .D(\register[11][3] ), .S0(n1472), .S1(n1431), .Y(
        n1162) );
  MXI4X1 U743 ( .A(\register[24][3] ), .B(\register[25][3] ), .C(
        \register[26][3] ), .D(\register[27][3] ), .S0(n1471), .S1(n1430), .Y(
        n1158) );
  MXI4X1 U744 ( .A(\register[8][1] ), .B(\register[9][1] ), .C(
        \register[10][1] ), .D(\register[11][1] ), .S0(n1470), .S1(n1429), .Y(
        n1146) );
  MXI4X1 U745 ( .A(\register[24][1] ), .B(\register[25][1] ), .C(
        \register[26][1] ), .D(\register[27][1] ), .S0(n1470), .S1(n1429), .Y(
        n1142) );
  MXI4X1 U746 ( .A(\register[8][0] ), .B(\register[9][0] ), .C(
        \register[10][0] ), .D(\register[11][0] ), .S0(n1470), .S1(n1429), .Y(
        n1138) );
  MXI4X1 U747 ( .A(\register[8][0] ), .B(\register[9][0] ), .C(
        \register[10][0] ), .D(\register[11][0] ), .S0(n1894), .S1(n1853), .Y(
        n1562) );
  MXI4X1 U748 ( .A(\register[24][1] ), .B(\register[25][1] ), .C(
        \register[26][1] ), .D(\register[27][1] ), .S0(n1894), .S1(n1853), .Y(
        n1566) );
  MXI4X1 U749 ( .A(\register[8][1] ), .B(\register[9][1] ), .C(
        \register[10][1] ), .D(\register[11][1] ), .S0(n1894), .S1(n1853), .Y(
        n1570) );
  MXI4X1 U750 ( .A(\register[24][2] ), .B(\register[25][2] ), .C(
        \register[26][2] ), .D(\register[27][2] ), .S0(n1895), .S1(n1854), .Y(
        n1574) );
  MXI4X1 U751 ( .A(\register[8][2] ), .B(\register[9][2] ), .C(
        \register[10][2] ), .D(\register[11][2] ), .S0(n1895), .S1(n1854), .Y(
        n1578) );
  MXI4X1 U752 ( .A(\register[24][3] ), .B(\register[25][3] ), .C(
        \register[26][3] ), .D(\register[27][3] ), .S0(n1895), .S1(n1854), .Y(
        n1582) );
  MXI4X1 U753 ( .A(\register[8][3] ), .B(\register[9][3] ), .C(
        \register[10][3] ), .D(\register[11][3] ), .S0(n1896), .S1(n1855), .Y(
        n1586) );
  MX4X1 U754 ( .A(n1204), .B(n1202), .C(n1203), .D(n1201), .S0(n1396), .S1(
        n1404), .Y(n17) );
  MX4X1 U755 ( .A(n1200), .B(n1198), .C(n1199), .D(n1197), .S0(n1396), .S1(
        n1404), .Y(n18) );
  MXI4X1 U756 ( .A(\register[0][8] ), .B(\register[1][8] ), .C(
        \register[2][8] ), .D(\register[3][8] ), .S0(n1475), .S1(n1434), .Y(
        n1204) );
  MXI2X1 U757 ( .A(n1501), .B(n1502), .S0(n1813), .Y(ReadData2_o[4]) );
  MX4X1 U758 ( .A(n1596), .B(n1594), .C(n1595), .D(n1593), .S0(n1819), .S1(
        n1827), .Y(n1501) );
  MX4X1 U759 ( .A(n1592), .B(n1590), .C(n1591), .D(n1589), .S0(n1819), .S1(
        n1827), .Y(n1502) );
  MXI4X1 U760 ( .A(\register[0][4] ), .B(\register[1][4] ), .C(
        \register[2][4] ), .D(\register[3][4] ), .S0(n1896), .S1(n1855), .Y(
        n1596) );
  MXI2X1 U761 ( .A(n1503), .B(n1504), .S0(n1813), .Y(ReadData2_o[5]) );
  MX4X1 U762 ( .A(n1604), .B(n1602), .C(n1603), .D(n1601), .S0(n1819), .S1(
        n1827), .Y(n1503) );
  MX4X1 U763 ( .A(n1600), .B(n1598), .C(n1599), .D(n1597), .S0(n1819), .S1(
        n1827), .Y(n1504) );
  MXI4X1 U764 ( .A(\register[0][5] ), .B(\register[1][5] ), .C(
        \register[2][5] ), .D(\register[3][5] ), .S0(n1897), .S1(n1856), .Y(
        n1604) );
  MX4X1 U765 ( .A(n1176), .B(n1174), .C(n1175), .D(n1173), .S0(n1395), .S1(
        n1403), .Y(n12) );
  MX4X1 U766 ( .A(n1180), .B(n1178), .C(n1179), .D(n1177), .S0(n1395), .S1(
        n1403), .Y(n11) );
  MXI4X1 U767 ( .A(\register[28][5] ), .B(\register[29][5] ), .C(
        \register[30][5] ), .D(\register[31][5] ), .S0(n1473), .S1(n1432), .Y(
        n1173) );
  MX4X1 U768 ( .A(n1168), .B(n1166), .C(n1167), .D(n1165), .S0(n1395), .S1(
        n1403), .Y(n10) );
  MX4X1 U769 ( .A(n1172), .B(n1170), .C(n1171), .D(n1169), .S0(n1395), .S1(
        n1403), .Y(n9) );
  MXI4X1 U770 ( .A(\register[28][4] ), .B(\register[29][4] ), .C(
        \register[30][4] ), .D(\register[31][4] ), .S0(n1472), .S1(n1431), .Y(
        n1165) );
  MX4X1 U771 ( .A(n1184), .B(n1182), .C(n1183), .D(n1181), .S0(n1395), .S1(
        n1404), .Y(n14) );
  MX4X1 U772 ( .A(n1188), .B(n1186), .C(n1187), .D(n1185), .S0(n1395), .S1(
        n1404), .Y(n13) );
  MXI4X1 U773 ( .A(\register[28][6] ), .B(\register[29][6] ), .C(
        \register[30][6] ), .D(\register[31][6] ), .S0(n1473), .S1(n1432), .Y(
        n1181) );
  MX4X1 U774 ( .A(n1192), .B(n1190), .C(n1191), .D(n1189), .S0(n1395), .S1(
        n1404), .Y(n16) );
  MX4X1 U775 ( .A(n1196), .B(n1194), .C(n1195), .D(n1193), .S0(n1395), .S1(
        n1404), .Y(n15) );
  MXI4X1 U776 ( .A(\register[24][7] ), .B(\register[25][7] ), .C(
        \register[26][7] ), .D(\register[27][7] ), .S0(n1474), .S1(n1433), .Y(
        n1190) );
  MXI2X1 U777 ( .A(n1505), .B(n1506), .S0(n1813), .Y(ReadData2_o[6]) );
  MX4X1 U778 ( .A(n1608), .B(n1606), .C(n1607), .D(n1605), .S0(n1819), .S1(
        n1828), .Y(n1506) );
  MX4X1 U779 ( .A(n1612), .B(n1610), .C(n1611), .D(n1609), .S0(n1819), .S1(
        n1828), .Y(n1505) );
  MXI4X1 U780 ( .A(\register[24][6] ), .B(\register[25][6] ), .C(
        \register[26][6] ), .D(\register[27][6] ), .S0(n1897), .S1(n1856), .Y(
        n1606) );
  MXI2X1 U781 ( .A(n1507), .B(n1508), .S0(n1813), .Y(ReadData2_o[7]) );
  MX4X1 U782 ( .A(n1616), .B(n1614), .C(n1615), .D(n1613), .S0(n1819), .S1(
        n1828), .Y(n1508) );
  MX4X1 U783 ( .A(n1620), .B(n1618), .C(n1619), .D(n1617), .S0(n1819), .S1(
        n1828), .Y(n1507) );
  MXI4X1 U784 ( .A(\register[28][7] ), .B(\register[29][7] ), .C(
        \register[30][7] ), .D(\register[31][7] ), .S0(n1898), .S1(n1857), .Y(
        n1613) );
  MXI2X1 U785 ( .A(n1509), .B(n1510), .S0(n1814), .Y(ReadData2_o[8]) );
  MX4X1 U786 ( .A(n1624), .B(n1622), .C(n1623), .D(n1621), .S0(n1820), .S1(
        n1828), .Y(n1510) );
  MX4X1 U787 ( .A(n1628), .B(n1626), .C(n1627), .D(n1625), .S0(n1820), .S1(
        n1828), .Y(n1509) );
  MXI4X1 U788 ( .A(\register[28][8] ), .B(\register[29][8] ), .C(
        \register[30][8] ), .D(\register[31][8] ), .S0(n1899), .S1(n1858), .Y(
        n1621) );
  MXI4X1 U789 ( .A(\register[4][5] ), .B(\register[5][5] ), .C(
        \register[6][5] ), .D(\register[7][5] ), .S0(n1473), .S1(n1432), .Y(
        n1179) );
  MXI4X1 U790 ( .A(\register[20][5] ), .B(\register[21][5] ), .C(
        \register[22][5] ), .D(\register[23][5] ), .S0(n1473), .S1(n1432), .Y(
        n1175) );
  MXI4X1 U791 ( .A(\register[20][8] ), .B(\register[21][8] ), .C(
        \register[22][8] ), .D(\register[23][8] ), .S0(n1475), .S1(n1434), .Y(
        n1199) );
  MXI4X1 U792 ( .A(\register[4][8] ), .B(\register[5][8] ), .C(
        \register[6][8] ), .D(\register[7][8] ), .S0(n1475), .S1(n1434), .Y(
        n1203) );
  MXI4X1 U793 ( .A(\register[4][4] ), .B(\register[5][4] ), .C(
        \register[6][4] ), .D(\register[7][4] ), .S0(n1472), .S1(n1431), .Y(
        n1171) );
  MXI4X1 U794 ( .A(\register[20][4] ), .B(\register[21][4] ), .C(
        \register[22][4] ), .D(\register[23][4] ), .S0(n1472), .S1(n1431), .Y(
        n1167) );
  MXI4X1 U795 ( .A(\register[4][6] ), .B(\register[5][6] ), .C(
        \register[6][6] ), .D(\register[7][6] ), .S0(n1474), .S1(n1433), .Y(
        n1187) );
  MXI4X1 U796 ( .A(\register[20][6] ), .B(\register[21][6] ), .C(
        \register[22][6] ), .D(\register[23][6] ), .S0(n1473), .S1(n1432), .Y(
        n1183) );
  MXI4X1 U797 ( .A(\register[4][7] ), .B(\register[5][7] ), .C(
        \register[6][7] ), .D(\register[7][7] ), .S0(n1474), .S1(n1433), .Y(
        n1195) );
  MXI4X1 U798 ( .A(\register[20][7] ), .B(\register[21][7] ), .C(
        \register[22][7] ), .D(\register[23][7] ), .S0(n1474), .S1(n1433), .Y(
        n1191) );
  MXI4X1 U799 ( .A(\register[20][4] ), .B(\register[21][4] ), .C(
        \register[22][4] ), .D(\register[23][4] ), .S0(n1896), .S1(n1855), .Y(
        n1591) );
  MXI4X1 U800 ( .A(\register[4][4] ), .B(\register[5][4] ), .C(
        \register[6][4] ), .D(\register[7][4] ), .S0(n1896), .S1(n1855), .Y(
        n1595) );
  MXI4X1 U801 ( .A(\register[20][5] ), .B(\register[21][5] ), .C(
        \register[22][5] ), .D(\register[23][5] ), .S0(n1897), .S1(n1856), .Y(
        n1599) );
  MXI4X1 U802 ( .A(\register[4][5] ), .B(\register[5][5] ), .C(
        \register[6][5] ), .D(\register[7][5] ), .S0(n1897), .S1(n1856), .Y(
        n1603) );
  MXI4X1 U803 ( .A(\register[4][6] ), .B(\register[5][6] ), .C(
        \register[6][6] ), .D(\register[7][6] ), .S0(n1898), .S1(n1857), .Y(
        n1611) );
  MXI4X1 U804 ( .A(\register[20][6] ), .B(\register[21][6] ), .C(
        \register[22][6] ), .D(\register[23][6] ), .S0(n1897), .S1(n1856), .Y(
        n1607) );
  MXI4X1 U805 ( .A(\register[4][7] ), .B(\register[5][7] ), .C(
        \register[6][7] ), .D(\register[7][7] ), .S0(n1898), .S1(n1857), .Y(
        n1619) );
  MXI4X1 U806 ( .A(\register[20][7] ), .B(\register[21][7] ), .C(
        \register[22][7] ), .D(\register[23][7] ), .S0(n1898), .S1(n1857), .Y(
        n1615) );
  MXI4X1 U807 ( .A(\register[4][8] ), .B(\register[5][8] ), .C(
        \register[6][8] ), .D(\register[7][8] ), .S0(n1899), .S1(n1858), .Y(
        n1627) );
  MXI4X1 U808 ( .A(\register[20][8] ), .B(\register[21][8] ), .C(
        \register[22][8] ), .D(\register[23][8] ), .S0(n1899), .S1(n1858), .Y(
        n1623) );
  MXI4X1 U809 ( .A(\register[0][5] ), .B(\register[1][5] ), .C(
        \register[2][5] ), .D(\register[3][5] ), .S0(n1473), .S1(n1432), .Y(
        n1180) );
  MXI4X1 U810 ( .A(\register[16][5] ), .B(\register[17][5] ), .C(
        \register[18][5] ), .D(\register[19][5] ), .S0(n1473), .S1(n1432), .Y(
        n1176) );
  MXI4X1 U811 ( .A(\register[16][8] ), .B(\register[17][8] ), .C(
        \register[18][8] ), .D(\register[19][8] ), .S0(n1475), .S1(n1434), .Y(
        n1200) );
  MXI4X1 U812 ( .A(\register[0][4] ), .B(\register[1][4] ), .C(
        \register[2][4] ), .D(\register[3][4] ), .S0(n1472), .S1(n1431), .Y(
        n1172) );
  MXI4X1 U813 ( .A(\register[16][4] ), .B(\register[17][4] ), .C(
        \register[18][4] ), .D(\register[19][4] ), .S0(n1472), .S1(n1431), .Y(
        n1168) );
  MXI4X1 U814 ( .A(\register[0][6] ), .B(\register[1][6] ), .C(
        \register[2][6] ), .D(\register[3][6] ), .S0(n1474), .S1(n1433), .Y(
        n1188) );
  MXI4X1 U815 ( .A(\register[16][6] ), .B(\register[17][6] ), .C(
        \register[18][6] ), .D(\register[19][6] ), .S0(n1473), .S1(n1432), .Y(
        n1184) );
  MXI4X1 U816 ( .A(\register[0][7] ), .B(\register[1][7] ), .C(
        \register[2][7] ), .D(\register[3][7] ), .S0(n1474), .S1(n1433), .Y(
        n1196) );
  MXI4X1 U817 ( .A(\register[16][7] ), .B(\register[17][7] ), .C(
        \register[18][7] ), .D(\register[19][7] ), .S0(n1474), .S1(n1433), .Y(
        n1192) );
  MXI4X1 U818 ( .A(\register[16][4] ), .B(\register[17][4] ), .C(
        \register[18][4] ), .D(\register[19][4] ), .S0(n1896), .S1(n1855), .Y(
        n1592) );
  MXI4X1 U819 ( .A(\register[16][5] ), .B(\register[17][5] ), .C(
        \register[18][5] ), .D(\register[19][5] ), .S0(n1897), .S1(n1856), .Y(
        n1600) );
  MXI4X1 U820 ( .A(\register[0][6] ), .B(\register[1][6] ), .C(
        \register[2][6] ), .D(\register[3][6] ), .S0(n1898), .S1(n1857), .Y(
        n1612) );
  MXI4X1 U821 ( .A(\register[16][6] ), .B(\register[17][6] ), .C(
        \register[18][6] ), .D(\register[19][6] ), .S0(n1897), .S1(n1856), .Y(
        n1608) );
  MXI4X1 U822 ( .A(\register[0][7] ), .B(\register[1][7] ), .C(
        \register[2][7] ), .D(\register[3][7] ), .S0(n1898), .S1(n1857), .Y(
        n1620) );
  MXI4X1 U823 ( .A(\register[16][7] ), .B(\register[17][7] ), .C(
        \register[18][7] ), .D(\register[19][7] ), .S0(n1898), .S1(n1857), .Y(
        n1616) );
  MXI4X1 U824 ( .A(\register[0][8] ), .B(\register[1][8] ), .C(
        \register[2][8] ), .D(\register[3][8] ), .S0(n1899), .S1(n1858), .Y(
        n1628) );
  MXI4X1 U825 ( .A(\register[16][8] ), .B(\register[17][8] ), .C(
        \register[18][8] ), .D(\register[19][8] ), .S0(n1899), .S1(n1858), .Y(
        n1624) );
  MXI4X1 U826 ( .A(\register[12][5] ), .B(\register[13][5] ), .C(
        \register[14][5] ), .D(\register[15][5] ), .S0(n1473), .S1(n1432), .Y(
        n1177) );
  MXI4X1 U827 ( .A(\register[28][8] ), .B(\register[29][8] ), .C(
        \register[30][8] ), .D(\register[31][8] ), .S0(n1475), .S1(n1434), .Y(
        n1197) );
  MXI4X1 U828 ( .A(\register[12][8] ), .B(\register[13][8] ), .C(
        \register[14][8] ), .D(\register[15][8] ), .S0(n1475), .S1(n1434), .Y(
        n1201) );
  MXI4X1 U829 ( .A(\register[12][4] ), .B(\register[13][4] ), .C(
        \register[14][4] ), .D(\register[15][4] ), .S0(n1472), .S1(n1431), .Y(
        n1169) );
  MXI4X1 U830 ( .A(\register[12][6] ), .B(\register[13][6] ), .C(
        \register[14][6] ), .D(\register[15][6] ), .S0(n1474), .S1(n1433), .Y(
        n1185) );
  MXI4X1 U831 ( .A(\register[12][7] ), .B(\register[13][7] ), .C(
        \register[14][7] ), .D(\register[15][7] ), .S0(n1474), .S1(n1433), .Y(
        n1193) );
  MXI4X1 U832 ( .A(\register[28][7] ), .B(\register[29][7] ), .C(
        \register[30][7] ), .D(\register[31][7] ), .S0(n1474), .S1(n1433), .Y(
        n1189) );
  MXI4X1 U833 ( .A(\register[28][4] ), .B(\register[29][4] ), .C(
        \register[30][4] ), .D(\register[31][4] ), .S0(n1896), .S1(n1855), .Y(
        n1589) );
  MXI4X1 U834 ( .A(\register[12][4] ), .B(\register[13][4] ), .C(
        \register[14][4] ), .D(\register[15][4] ), .S0(n1896), .S1(n1855), .Y(
        n1593) );
  MXI4X1 U835 ( .A(\register[28][5] ), .B(\register[29][5] ), .C(
        \register[30][5] ), .D(\register[31][5] ), .S0(n1897), .S1(n1856), .Y(
        n1597) );
  MXI4X1 U836 ( .A(\register[12][5] ), .B(\register[13][5] ), .C(
        \register[14][5] ), .D(\register[15][5] ), .S0(n1897), .S1(n1856), .Y(
        n1601) );
  MXI4X1 U837 ( .A(\register[12][6] ), .B(\register[13][6] ), .C(
        \register[14][6] ), .D(\register[15][6] ), .S0(n1898), .S1(n1857), .Y(
        n1609) );
  MXI4X1 U838 ( .A(\register[28][6] ), .B(\register[29][6] ), .C(
        \register[30][6] ), .D(\register[31][6] ), .S0(n1897), .S1(n1856), .Y(
        n1605) );
  MXI4X1 U839 ( .A(\register[12][7] ), .B(\register[13][7] ), .C(
        \register[14][7] ), .D(\register[15][7] ), .S0(n1898), .S1(n1857), .Y(
        n1617) );
  MXI4X1 U840 ( .A(\register[12][8] ), .B(\register[13][8] ), .C(
        \register[14][8] ), .D(\register[15][8] ), .S0(n1899), .S1(n1858), .Y(
        n1625) );
  MXI4X1 U841 ( .A(\register[8][5] ), .B(\register[9][5] ), .C(
        \register[10][5] ), .D(\register[11][5] ), .S0(n1473), .S1(n1432), .Y(
        n1178) );
  MXI4X1 U842 ( .A(\register[24][5] ), .B(\register[25][5] ), .C(
        \register[26][5] ), .D(\register[27][5] ), .S0(n1473), .S1(n1432), .Y(
        n1174) );
  MXI4X1 U843 ( .A(\register[24][8] ), .B(\register[25][8] ), .C(
        \register[26][8] ), .D(\register[27][8] ), .S0(n1475), .S1(n1434), .Y(
        n1198) );
  MXI4X1 U844 ( .A(\register[8][8] ), .B(\register[9][8] ), .C(
        \register[10][8] ), .D(\register[11][8] ), .S0(n1475), .S1(n1434), .Y(
        n1202) );
  MXI4X1 U845 ( .A(\register[8][4] ), .B(\register[9][4] ), .C(
        \register[10][4] ), .D(\register[11][4] ), .S0(n1472), .S1(n1431), .Y(
        n1170) );
  MXI4X1 U846 ( .A(\register[24][4] ), .B(\register[25][4] ), .C(
        \register[26][4] ), .D(\register[27][4] ), .S0(n1472), .S1(n1431), .Y(
        n1166) );
  MXI4X1 U847 ( .A(\register[8][6] ), .B(\register[9][6] ), .C(
        \register[10][6] ), .D(\register[11][6] ), .S0(n1474), .S1(n1433), .Y(
        n1186) );
  MXI4X1 U848 ( .A(\register[24][6] ), .B(\register[25][6] ), .C(
        \register[26][6] ), .D(\register[27][6] ), .S0(n1473), .S1(n1432), .Y(
        n1182) );
  MXI4X1 U849 ( .A(\register[8][7] ), .B(\register[9][7] ), .C(
        \register[10][7] ), .D(\register[11][7] ), .S0(n1474), .S1(n1433), .Y(
        n1194) );
  MXI4X1 U850 ( .A(\register[24][4] ), .B(\register[25][4] ), .C(
        \register[26][4] ), .D(\register[27][4] ), .S0(n1896), .S1(n1855), .Y(
        n1590) );
  MXI4X1 U851 ( .A(\register[8][4] ), .B(\register[9][4] ), .C(
        \register[10][4] ), .D(\register[11][4] ), .S0(n1896), .S1(n1855), .Y(
        n1594) );
  MXI4X1 U852 ( .A(\register[24][5] ), .B(\register[25][5] ), .C(
        \register[26][5] ), .D(\register[27][5] ), .S0(n1897), .S1(n1856), .Y(
        n1598) );
  MXI4X1 U853 ( .A(\register[8][5] ), .B(\register[9][5] ), .C(
        \register[10][5] ), .D(\register[11][5] ), .S0(n1897), .S1(n1856), .Y(
        n1602) );
  MXI4X1 U854 ( .A(\register[8][6] ), .B(\register[9][6] ), .C(
        \register[10][6] ), .D(\register[11][6] ), .S0(n1898), .S1(n1857), .Y(
        n1610) );
  MXI4X1 U855 ( .A(\register[8][7] ), .B(\register[9][7] ), .C(
        \register[10][7] ), .D(\register[11][7] ), .S0(n1898), .S1(n1857), .Y(
        n1618) );
  MXI4X1 U856 ( .A(\register[24][7] ), .B(\register[25][7] ), .C(
        \register[26][7] ), .D(\register[27][7] ), .S0(n1898), .S1(n1857), .Y(
        n1614) );
  MXI4X1 U857 ( .A(\register[8][8] ), .B(\register[9][8] ), .C(
        \register[10][8] ), .D(\register[11][8] ), .S0(n1899), .S1(n1858), .Y(
        n1626) );
  MXI4X1 U858 ( .A(\register[24][8] ), .B(\register[25][8] ), .C(
        \register[26][8] ), .D(\register[27][8] ), .S0(n1899), .S1(n1858), .Y(
        n1622) );
  OAI2BB2XL U859 ( .B0(n2012), .B1(n2266), .A0N(\register[30][0] ), .A1N(n2268), .Y(n114) );
  OAI2BB2XL U860 ( .B0(n2009), .B1(n2266), .A0N(\register[30][1] ), .A1N(n2269), .Y(n115) );
  OAI2BB2XL U861 ( .B0(n2006), .B1(n2266), .A0N(\register[30][2] ), .A1N(n2269), .Y(n116) );
  OAI2BB2XL U862 ( .B0(n2003), .B1(n2266), .A0N(\register[30][3] ), .A1N(n2269), .Y(n117) );
  OAI2BB2XL U863 ( .B0(n2000), .B1(n2266), .A0N(\register[30][4] ), .A1N(n2269), .Y(n118) );
  OAI2BB2XL U864 ( .B0(n1997), .B1(n2266), .A0N(\register[30][5] ), .A1N(n2269), .Y(n119) );
  OAI2BB2XL U865 ( .B0(n1994), .B1(n2266), .A0N(\register[30][6] ), .A1N(n2269), .Y(n120) );
  OAI2BB2XL U866 ( .B0(n1991), .B1(n2266), .A0N(\register[30][7] ), .A1N(n2269), .Y(n121) );
  OAI2BB2XL U867 ( .B0(n1988), .B1(n2267), .A0N(\register[30][8] ), .A1N(n2269), .Y(n122) );
  OAI2BB2XL U868 ( .B0(n1985), .B1(n2267), .A0N(\register[30][9] ), .A1N(n2269), .Y(n123) );
  OAI2BB2XL U869 ( .B0(n1982), .B1(n2267), .A0N(\register[30][10] ), .A1N(
        n2269), .Y(n124) );
  OAI2BB2XL U870 ( .B0(n1979), .B1(n2267), .A0N(\register[30][11] ), .A1N(
        n2269), .Y(n125) );
  OAI2BB2XL U871 ( .B0(n1976), .B1(n2267), .A0N(\register[30][12] ), .A1N(
        n2269), .Y(n126) );
  OAI2BB2XL U872 ( .B0(n1973), .B1(n2267), .A0N(\register[30][13] ), .A1N(
        n2269), .Y(n127) );
  OAI2BB2XL U873 ( .B0(n1970), .B1(n2267), .A0N(\register[30][14] ), .A1N(
        n2269), .Y(n128) );
  OAI2BB2XL U874 ( .B0(n1967), .B1(n2267), .A0N(\register[30][15] ), .A1N(
        n2269), .Y(n129) );
  OAI2BB2XL U875 ( .B0(n1964), .B1(n2268), .A0N(\register[30][16] ), .A1N(
        n2269), .Y(n130) );
  OAI2BB2XL U876 ( .B0(n1961), .B1(n2268), .A0N(\register[30][17] ), .A1N(
        n2269), .Y(n131) );
  OAI2BB2XL U877 ( .B0(n1958), .B1(n2267), .A0N(\register[30][18] ), .A1N(
        n2269), .Y(n132) );
  OAI2BB2XL U878 ( .B0(n1955), .B1(n2268), .A0N(\register[30][19] ), .A1N(
        n2269), .Y(n133) );
  OAI2BB2XL U879 ( .B0(n1952), .B1(n2268), .A0N(\register[30][20] ), .A1N(
        n2269), .Y(n134) );
  OAI2BB2XL U880 ( .B0(n1949), .B1(n2268), .A0N(\register[30][21] ), .A1N(
        n2268), .Y(n135) );
  OAI2BB2XL U881 ( .B0(n1946), .B1(n2268), .A0N(\register[30][22] ), .A1N(
        n2268), .Y(n136) );
  OAI2BB2XL U882 ( .B0(n1943), .B1(n2268), .A0N(\register[30][23] ), .A1N(
        n2268), .Y(n137) );
  OAI2BB2XL U883 ( .B0(n1940), .B1(n2268), .A0N(\register[30][24] ), .A1N(
        n2268), .Y(n138) );
  OAI2BB2XL U884 ( .B0(n1937), .B1(n2267), .A0N(\register[30][25] ), .A1N(
        n2268), .Y(n139) );
  OAI2BB2XL U885 ( .B0(n1934), .B1(n2267), .A0N(\register[30][26] ), .A1N(
        n2268), .Y(n140) );
  OAI2BB2XL U886 ( .B0(n1931), .B1(n2267), .A0N(\register[30][27] ), .A1N(
        n2268), .Y(n141) );
  OAI2BB2XL U887 ( .B0(n1928), .B1(n2266), .A0N(\register[30][28] ), .A1N(
        n2268), .Y(n142) );
  OAI2BB2XL U888 ( .B0(n1925), .B1(n2266), .A0N(\register[30][29] ), .A1N(
        n2268), .Y(n143) );
  OAI2BB2XL U889 ( .B0(n1922), .B1(n2266), .A0N(\register[30][30] ), .A1N(
        n2268), .Y(n144) );
  OAI2BB2XL U890 ( .B0(n1919), .B1(n2266), .A0N(\register[30][31] ), .A1N(
        n2268), .Y(n145) );
  OAI2BB2XL U891 ( .B0(n2012), .B1(n2262), .A0N(\register[29][0] ), .A1N(n2264), .Y(n146) );
  OAI2BB2XL U892 ( .B0(n2009), .B1(n2262), .A0N(\register[29][1] ), .A1N(n2265), .Y(n147) );
  OAI2BB2XL U893 ( .B0(n2006), .B1(n2262), .A0N(\register[29][2] ), .A1N(n2265), .Y(n148) );
  OAI2BB2XL U894 ( .B0(n2003), .B1(n2262), .A0N(\register[29][3] ), .A1N(n2265), .Y(n149) );
  OAI2BB2XL U895 ( .B0(n2000), .B1(n2262), .A0N(\register[29][4] ), .A1N(n2265), .Y(n150) );
  OAI2BB2XL U896 ( .B0(n1997), .B1(n2262), .A0N(\register[29][5] ), .A1N(n2265), .Y(n151) );
  OAI2BB2XL U897 ( .B0(n1994), .B1(n2262), .A0N(\register[29][6] ), .A1N(n2265), .Y(n152) );
  OAI2BB2XL U898 ( .B0(n1991), .B1(n2262), .A0N(\register[29][7] ), .A1N(n2265), .Y(n153) );
  OAI2BB2XL U899 ( .B0(n1988), .B1(n2263), .A0N(\register[29][8] ), .A1N(n2265), .Y(n154) );
  OAI2BB2XL U900 ( .B0(n1985), .B1(n2263), .A0N(\register[29][9] ), .A1N(n2265), .Y(n155) );
  OAI2BB2XL U901 ( .B0(n1982), .B1(n2263), .A0N(\register[29][10] ), .A1N(
        n2265), .Y(n156) );
  OAI2BB2XL U902 ( .B0(n1979), .B1(n2263), .A0N(\register[29][11] ), .A1N(
        n2265), .Y(n157) );
  OAI2BB2XL U903 ( .B0(n1976), .B1(n2263), .A0N(\register[29][12] ), .A1N(
        n2265), .Y(n158) );
  OAI2BB2XL U904 ( .B0(n1973), .B1(n2263), .A0N(\register[29][13] ), .A1N(
        n2265), .Y(n159) );
  OAI2BB2XL U905 ( .B0(n1970), .B1(n2263), .A0N(\register[29][14] ), .A1N(
        n2265), .Y(n160) );
  OAI2BB2XL U906 ( .B0(n1967), .B1(n2263), .A0N(\register[29][15] ), .A1N(
        n2265), .Y(n161) );
  OAI2BB2XL U907 ( .B0(n1964), .B1(n2264), .A0N(\register[29][16] ), .A1N(
        n2265), .Y(n162) );
  OAI2BB2XL U908 ( .B0(n1961), .B1(n2264), .A0N(\register[29][17] ), .A1N(
        n2265), .Y(n163) );
  OAI2BB2XL U909 ( .B0(n1958), .B1(n2263), .A0N(\register[29][18] ), .A1N(
        n2265), .Y(n164) );
  OAI2BB2XL U910 ( .B0(n1955), .B1(n2264), .A0N(\register[29][19] ), .A1N(
        n2265), .Y(n165) );
  OAI2BB2XL U911 ( .B0(n1952), .B1(n2264), .A0N(\register[29][20] ), .A1N(
        n2265), .Y(n166) );
  OAI2BB2XL U912 ( .B0(n1949), .B1(n2264), .A0N(\register[29][21] ), .A1N(
        n2264), .Y(n167) );
  OAI2BB2XL U913 ( .B0(n1946), .B1(n2264), .A0N(\register[29][22] ), .A1N(
        n2264), .Y(n168) );
  OAI2BB2XL U914 ( .B0(n1943), .B1(n2264), .A0N(\register[29][23] ), .A1N(
        n2264), .Y(n169) );
  OAI2BB2XL U915 ( .B0(n1940), .B1(n2264), .A0N(\register[29][24] ), .A1N(
        n2264), .Y(n170) );
  OAI2BB2XL U916 ( .B0(n1937), .B1(n2263), .A0N(\register[29][25] ), .A1N(
        n2264), .Y(n171) );
  OAI2BB2XL U917 ( .B0(n1934), .B1(n2263), .A0N(\register[29][26] ), .A1N(
        n2264), .Y(n172) );
  OAI2BB2XL U918 ( .B0(n1931), .B1(n2263), .A0N(\register[29][27] ), .A1N(
        n2264), .Y(n173) );
  OAI2BB2XL U919 ( .B0(n1928), .B1(n2262), .A0N(\register[29][28] ), .A1N(
        n2264), .Y(n174) );
  OAI2BB2XL U920 ( .B0(n1925), .B1(n2262), .A0N(\register[29][29] ), .A1N(
        n2264), .Y(n175) );
  OAI2BB2XL U921 ( .B0(n1922), .B1(n2262), .A0N(\register[29][30] ), .A1N(
        n2264), .Y(n176) );
  OAI2BB2XL U922 ( .B0(n1919), .B1(n2262), .A0N(\register[29][31] ), .A1N(
        n2264), .Y(n177) );
  OAI2BB2XL U923 ( .B0(n2012), .B1(n2258), .A0N(\register[28][0] ), .A1N(n2260), .Y(n178) );
  OAI2BB2XL U924 ( .B0(n2009), .B1(n2258), .A0N(\register[28][1] ), .A1N(n2261), .Y(n179) );
  OAI2BB2XL U925 ( .B0(n2006), .B1(n2258), .A0N(\register[28][2] ), .A1N(n2261), .Y(n180) );
  OAI2BB2XL U926 ( .B0(n2003), .B1(n2258), .A0N(\register[28][3] ), .A1N(n2261), .Y(n181) );
  OAI2BB2XL U927 ( .B0(n2000), .B1(n2258), .A0N(\register[28][4] ), .A1N(n2261), .Y(n182) );
  OAI2BB2XL U928 ( .B0(n1997), .B1(n2258), .A0N(\register[28][5] ), .A1N(n2261), .Y(n183) );
  OAI2BB2XL U929 ( .B0(n1994), .B1(n2258), .A0N(\register[28][6] ), .A1N(n2261), .Y(n184) );
  OAI2BB2XL U930 ( .B0(n1991), .B1(n2258), .A0N(\register[28][7] ), .A1N(n2261), .Y(n185) );
  OAI2BB2XL U931 ( .B0(n1988), .B1(n2259), .A0N(\register[28][8] ), .A1N(n2261), .Y(n186) );
  OAI2BB2XL U932 ( .B0(n1985), .B1(n2259), .A0N(\register[28][9] ), .A1N(n2261), .Y(n187) );
  OAI2BB2XL U933 ( .B0(n1982), .B1(n2259), .A0N(\register[28][10] ), .A1N(
        n2261), .Y(n188) );
  OAI2BB2XL U934 ( .B0(n1979), .B1(n2259), .A0N(\register[28][11] ), .A1N(
        n2261), .Y(n189) );
  OAI2BB2XL U935 ( .B0(n1976), .B1(n2259), .A0N(\register[28][12] ), .A1N(
        n2261), .Y(n190) );
  OAI2BB2XL U936 ( .B0(n1973), .B1(n2259), .A0N(\register[28][13] ), .A1N(
        n2261), .Y(n191) );
  OAI2BB2XL U937 ( .B0(n1970), .B1(n2259), .A0N(\register[28][14] ), .A1N(
        n2261), .Y(n192) );
  OAI2BB2XL U938 ( .B0(n1967), .B1(n2259), .A0N(\register[28][15] ), .A1N(
        n2261), .Y(n193) );
  OAI2BB2XL U939 ( .B0(n1964), .B1(n2260), .A0N(\register[28][16] ), .A1N(
        n2261), .Y(n194) );
  OAI2BB2XL U940 ( .B0(n1961), .B1(n2260), .A0N(\register[28][17] ), .A1N(
        n2261), .Y(n195) );
  OAI2BB2XL U941 ( .B0(n1958), .B1(n2259), .A0N(\register[28][18] ), .A1N(
        n2261), .Y(n196) );
  OAI2BB2XL U942 ( .B0(n1955), .B1(n2260), .A0N(\register[28][19] ), .A1N(
        n2261), .Y(n197) );
  OAI2BB2XL U943 ( .B0(n1952), .B1(n2260), .A0N(\register[28][20] ), .A1N(
        n2261), .Y(n198) );
  OAI2BB2XL U944 ( .B0(n1949), .B1(n2260), .A0N(\register[28][21] ), .A1N(
        n2260), .Y(n199) );
  OAI2BB2XL U945 ( .B0(n1946), .B1(n2260), .A0N(\register[28][22] ), .A1N(
        n2260), .Y(n200) );
  OAI2BB2XL U946 ( .B0(n1943), .B1(n2260), .A0N(\register[28][23] ), .A1N(
        n2260), .Y(n201) );
  OAI2BB2XL U947 ( .B0(n1940), .B1(n2260), .A0N(\register[28][24] ), .A1N(
        n2260), .Y(n202) );
  OAI2BB2XL U948 ( .B0(n1937), .B1(n2259), .A0N(\register[28][25] ), .A1N(
        n2260), .Y(n203) );
  OAI2BB2XL U949 ( .B0(n1934), .B1(n2259), .A0N(\register[28][26] ), .A1N(
        n2260), .Y(n204) );
  OAI2BB2XL U950 ( .B0(n1931), .B1(n2259), .A0N(\register[28][27] ), .A1N(
        n2260), .Y(n205) );
  OAI2BB2XL U951 ( .B0(n1928), .B1(n2258), .A0N(\register[28][28] ), .A1N(
        n2260), .Y(n206) );
  OAI2BB2XL U952 ( .B0(n1925), .B1(n2258), .A0N(\register[28][29] ), .A1N(
        n2260), .Y(n207) );
  OAI2BB2XL U953 ( .B0(n1922), .B1(n2258), .A0N(\register[28][30] ), .A1N(
        n2260), .Y(n208) );
  OAI2BB2XL U954 ( .B0(n1919), .B1(n2258), .A0N(\register[28][31] ), .A1N(
        n2260), .Y(n209) );
  OAI2BB2XL U955 ( .B0(n2012), .B1(n2254), .A0N(\register[27][0] ), .A1N(n2256), .Y(n210) );
  OAI2BB2XL U956 ( .B0(n2009), .B1(n2254), .A0N(\register[27][1] ), .A1N(n2257), .Y(n211) );
  OAI2BB2XL U957 ( .B0(n2006), .B1(n2254), .A0N(\register[27][2] ), .A1N(n2257), .Y(n212) );
  OAI2BB2XL U958 ( .B0(n2003), .B1(n2254), .A0N(\register[27][3] ), .A1N(n2257), .Y(n213) );
  OAI2BB2XL U959 ( .B0(n2000), .B1(n2254), .A0N(\register[27][4] ), .A1N(n2257), .Y(n214) );
  OAI2BB2XL U960 ( .B0(n1997), .B1(n2254), .A0N(\register[27][5] ), .A1N(n2257), .Y(n215) );
  OAI2BB2XL U961 ( .B0(n1994), .B1(n2254), .A0N(\register[27][6] ), .A1N(n2257), .Y(n216) );
  OAI2BB2XL U962 ( .B0(n1991), .B1(n2254), .A0N(\register[27][7] ), .A1N(n2257), .Y(n217) );
  OAI2BB2XL U963 ( .B0(n1988), .B1(n2255), .A0N(\register[27][8] ), .A1N(n2257), .Y(n218) );
  OAI2BB2XL U964 ( .B0(n1985), .B1(n2255), .A0N(\register[27][9] ), .A1N(n2257), .Y(n219) );
  OAI2BB2XL U965 ( .B0(n1982), .B1(n2255), .A0N(\register[27][10] ), .A1N(
        n2257), .Y(n220) );
  OAI2BB2XL U966 ( .B0(n1979), .B1(n2255), .A0N(\register[27][11] ), .A1N(
        n2257), .Y(n221) );
  OAI2BB2XL U967 ( .B0(n1976), .B1(n2255), .A0N(\register[27][12] ), .A1N(
        n2257), .Y(n222) );
  OAI2BB2XL U968 ( .B0(n1973), .B1(n2255), .A0N(\register[27][13] ), .A1N(
        n2257), .Y(n223) );
  OAI2BB2XL U969 ( .B0(n1970), .B1(n2255), .A0N(\register[27][14] ), .A1N(
        n2257), .Y(n224) );
  OAI2BB2XL U970 ( .B0(n1967), .B1(n2255), .A0N(\register[27][15] ), .A1N(
        n2257), .Y(n225) );
  OAI2BB2XL U971 ( .B0(n1964), .B1(n2256), .A0N(\register[27][16] ), .A1N(
        n2257), .Y(n226) );
  OAI2BB2XL U972 ( .B0(n1961), .B1(n2256), .A0N(\register[27][17] ), .A1N(
        n2257), .Y(n227) );
  OAI2BB2XL U973 ( .B0(n1958), .B1(n2255), .A0N(\register[27][18] ), .A1N(
        n2257), .Y(n228) );
  OAI2BB2XL U974 ( .B0(n1955), .B1(n2256), .A0N(\register[27][19] ), .A1N(
        n2257), .Y(n229) );
  OAI2BB2XL U975 ( .B0(n1952), .B1(n2256), .A0N(\register[27][20] ), .A1N(
        n2257), .Y(n230) );
  OAI2BB2XL U976 ( .B0(n1949), .B1(n2256), .A0N(\register[27][21] ), .A1N(
        n2256), .Y(n231) );
  OAI2BB2XL U977 ( .B0(n1946), .B1(n2256), .A0N(\register[27][22] ), .A1N(
        n2256), .Y(n232) );
  OAI2BB2XL U978 ( .B0(n1943), .B1(n2256), .A0N(\register[27][23] ), .A1N(
        n2256), .Y(n233) );
  OAI2BB2XL U979 ( .B0(n1940), .B1(n2256), .A0N(\register[27][24] ), .A1N(
        n2256), .Y(n234) );
  OAI2BB2XL U980 ( .B0(n1937), .B1(n2255), .A0N(\register[27][25] ), .A1N(
        n2256), .Y(n235) );
  OAI2BB2XL U981 ( .B0(n1934), .B1(n2255), .A0N(\register[27][26] ), .A1N(
        n2256), .Y(n236) );
  OAI2BB2XL U982 ( .B0(n1931), .B1(n2255), .A0N(\register[27][27] ), .A1N(
        n2256), .Y(n237) );
  OAI2BB2XL U983 ( .B0(n1928), .B1(n2254), .A0N(\register[27][28] ), .A1N(
        n2256), .Y(n238) );
  OAI2BB2XL U984 ( .B0(n1925), .B1(n2254), .A0N(\register[27][29] ), .A1N(
        n2256), .Y(n239) );
  OAI2BB2XL U985 ( .B0(n1922), .B1(n2254), .A0N(\register[27][30] ), .A1N(
        n2256), .Y(n240) );
  OAI2BB2XL U986 ( .B0(n1919), .B1(n2254), .A0N(\register[27][31] ), .A1N(
        n2256), .Y(n241) );
  OAI2BB2XL U987 ( .B0(n2012), .B1(n2250), .A0N(\register[26][0] ), .A1N(n2252), .Y(n242) );
  OAI2BB2XL U988 ( .B0(n2009), .B1(n2250), .A0N(\register[26][1] ), .A1N(n2253), .Y(n243) );
  OAI2BB2XL U989 ( .B0(n2006), .B1(n2250), .A0N(\register[26][2] ), .A1N(n2253), .Y(n244) );
  OAI2BB2XL U990 ( .B0(n2003), .B1(n2250), .A0N(\register[26][3] ), .A1N(n2253), .Y(n245) );
  OAI2BB2XL U991 ( .B0(n2000), .B1(n2250), .A0N(\register[26][4] ), .A1N(n2253), .Y(n246) );
  OAI2BB2XL U992 ( .B0(n1997), .B1(n2250), .A0N(\register[26][5] ), .A1N(n2253), .Y(n247) );
  OAI2BB2XL U993 ( .B0(n1994), .B1(n2250), .A0N(\register[26][6] ), .A1N(n2253), .Y(n248) );
  OAI2BB2XL U994 ( .B0(n1991), .B1(n2250), .A0N(\register[26][7] ), .A1N(n2253), .Y(n249) );
  OAI2BB2XL U995 ( .B0(n1988), .B1(n2251), .A0N(\register[26][8] ), .A1N(n2253), .Y(n250) );
  OAI2BB2XL U996 ( .B0(n1985), .B1(n2251), .A0N(\register[26][9] ), .A1N(n2253), .Y(n251) );
  OAI2BB2XL U997 ( .B0(n1982), .B1(n2251), .A0N(\register[26][10] ), .A1N(
        n2253), .Y(n252) );
  OAI2BB2XL U998 ( .B0(n1979), .B1(n2251), .A0N(\register[26][11] ), .A1N(
        n2253), .Y(n253) );
  OAI2BB2XL U999 ( .B0(n1976), .B1(n2251), .A0N(\register[26][12] ), .A1N(
        n2253), .Y(n254) );
  OAI2BB2XL U1000 ( .B0(n1973), .B1(n2251), .A0N(\register[26][13] ), .A1N(
        n2253), .Y(n255) );
  OAI2BB2XL U1001 ( .B0(n1970), .B1(n2251), .A0N(\register[26][14] ), .A1N(
        n2253), .Y(n256) );
  OAI2BB2XL U1002 ( .B0(n1967), .B1(n2251), .A0N(\register[26][15] ), .A1N(
        n2253), .Y(n257) );
  OAI2BB2XL U1003 ( .B0(n1964), .B1(n2252), .A0N(\register[26][16] ), .A1N(
        n2253), .Y(n258) );
  OAI2BB2XL U1004 ( .B0(n1961), .B1(n2252), .A0N(\register[26][17] ), .A1N(
        n2253), .Y(n259) );
  OAI2BB2XL U1005 ( .B0(n1958), .B1(n2251), .A0N(\register[26][18] ), .A1N(
        n2253), .Y(n260) );
  OAI2BB2XL U1006 ( .B0(n1955), .B1(n2252), .A0N(\register[26][19] ), .A1N(
        n2253), .Y(n261) );
  OAI2BB2XL U1007 ( .B0(n1952), .B1(n2252), .A0N(\register[26][20] ), .A1N(
        n2253), .Y(n262) );
  OAI2BB2XL U1008 ( .B0(n1949), .B1(n2252), .A0N(\register[26][21] ), .A1N(
        n2252), .Y(n263) );
  OAI2BB2XL U1009 ( .B0(n1946), .B1(n2252), .A0N(\register[26][22] ), .A1N(
        n2252), .Y(n264) );
  OAI2BB2XL U1010 ( .B0(n1943), .B1(n2252), .A0N(\register[26][23] ), .A1N(
        n2252), .Y(n265) );
  OAI2BB2XL U1011 ( .B0(n1940), .B1(n2252), .A0N(\register[26][24] ), .A1N(
        n2252), .Y(n266) );
  OAI2BB2XL U1012 ( .B0(n1937), .B1(n2251), .A0N(\register[26][25] ), .A1N(
        n2252), .Y(n267) );
  OAI2BB2XL U1013 ( .B0(n1934), .B1(n2251), .A0N(\register[26][26] ), .A1N(
        n2252), .Y(n268) );
  OAI2BB2XL U1014 ( .B0(n1931), .B1(n2251), .A0N(\register[26][27] ), .A1N(
        n2252), .Y(n269) );
  OAI2BB2XL U1015 ( .B0(n1928), .B1(n2250), .A0N(\register[26][28] ), .A1N(
        n2252), .Y(n270) );
  OAI2BB2XL U1016 ( .B0(n1925), .B1(n2250), .A0N(\register[26][29] ), .A1N(
        n2252), .Y(n271) );
  OAI2BB2XL U1017 ( .B0(n1922), .B1(n2250), .A0N(\register[26][30] ), .A1N(
        n2252), .Y(n272) );
  OAI2BB2XL U1018 ( .B0(n1919), .B1(n2250), .A0N(\register[26][31] ), .A1N(
        n2252), .Y(n273) );
  OAI2BB2XL U1019 ( .B0(n2012), .B1(n2246), .A0N(\register[25][0] ), .A1N(
        n2248), .Y(n274) );
  OAI2BB2XL U1020 ( .B0(n2009), .B1(n2246), .A0N(\register[25][1] ), .A1N(
        n2249), .Y(n275) );
  OAI2BB2XL U1021 ( .B0(n2006), .B1(n2246), .A0N(\register[25][2] ), .A1N(
        n2249), .Y(n276) );
  OAI2BB2XL U1022 ( .B0(n2003), .B1(n2246), .A0N(\register[25][3] ), .A1N(
        n2249), .Y(n277) );
  OAI2BB2XL U1023 ( .B0(n2000), .B1(n2246), .A0N(\register[25][4] ), .A1N(
        n2249), .Y(n278) );
  OAI2BB2XL U1024 ( .B0(n1997), .B1(n2246), .A0N(\register[25][5] ), .A1N(
        n2249), .Y(n279) );
  OAI2BB2XL U1025 ( .B0(n1994), .B1(n2246), .A0N(\register[25][6] ), .A1N(
        n2249), .Y(n280) );
  OAI2BB2XL U1026 ( .B0(n1991), .B1(n2246), .A0N(\register[25][7] ), .A1N(
        n2249), .Y(n281) );
  OAI2BB2XL U1027 ( .B0(n1988), .B1(n2247), .A0N(\register[25][8] ), .A1N(
        n2249), .Y(n282) );
  OAI2BB2XL U1028 ( .B0(n1985), .B1(n2247), .A0N(\register[25][9] ), .A1N(
        n2249), .Y(n283) );
  OAI2BB2XL U1029 ( .B0(n1982), .B1(n2247), .A0N(\register[25][10] ), .A1N(
        n2249), .Y(n284) );
  OAI2BB2XL U1030 ( .B0(n1979), .B1(n2247), .A0N(\register[25][11] ), .A1N(
        n2249), .Y(n285) );
  OAI2BB2XL U1031 ( .B0(n1976), .B1(n2247), .A0N(\register[25][12] ), .A1N(
        n2249), .Y(n286) );
  OAI2BB2XL U1032 ( .B0(n1973), .B1(n2247), .A0N(\register[25][13] ), .A1N(
        n2249), .Y(n287) );
  OAI2BB2XL U1033 ( .B0(n1970), .B1(n2247), .A0N(\register[25][14] ), .A1N(
        n2249), .Y(n288) );
  OAI2BB2XL U1034 ( .B0(n1967), .B1(n2247), .A0N(\register[25][15] ), .A1N(
        n2249), .Y(n289) );
  OAI2BB2XL U1035 ( .B0(n1964), .B1(n2248), .A0N(\register[25][16] ), .A1N(
        n2249), .Y(n290) );
  OAI2BB2XL U1036 ( .B0(n1961), .B1(n2248), .A0N(\register[25][17] ), .A1N(
        n2249), .Y(n291) );
  OAI2BB2XL U1037 ( .B0(n1958), .B1(n2247), .A0N(\register[25][18] ), .A1N(
        n2249), .Y(n292) );
  OAI2BB2XL U1038 ( .B0(n1955), .B1(n2248), .A0N(\register[25][19] ), .A1N(
        n2249), .Y(n293) );
  OAI2BB2XL U1039 ( .B0(n1952), .B1(n2248), .A0N(\register[25][20] ), .A1N(
        n2249), .Y(n294) );
  OAI2BB2XL U1040 ( .B0(n1949), .B1(n2248), .A0N(\register[25][21] ), .A1N(
        n2248), .Y(n295) );
  OAI2BB2XL U1041 ( .B0(n1946), .B1(n2248), .A0N(\register[25][22] ), .A1N(
        n2248), .Y(n296) );
  OAI2BB2XL U1042 ( .B0(n1943), .B1(n2248), .A0N(\register[25][23] ), .A1N(
        n2248), .Y(n297) );
  OAI2BB2XL U1043 ( .B0(n1940), .B1(n2248), .A0N(\register[25][24] ), .A1N(
        n2248), .Y(n298) );
  OAI2BB2XL U1044 ( .B0(n1937), .B1(n2247), .A0N(\register[25][25] ), .A1N(
        n2248), .Y(n299) );
  OAI2BB2XL U1045 ( .B0(n1934), .B1(n2247), .A0N(\register[25][26] ), .A1N(
        n2248), .Y(n300) );
  OAI2BB2XL U1046 ( .B0(n1931), .B1(n2247), .A0N(\register[25][27] ), .A1N(
        n2248), .Y(n301) );
  OAI2BB2XL U1047 ( .B0(n1928), .B1(n2246), .A0N(\register[25][28] ), .A1N(
        n2248), .Y(n302) );
  OAI2BB2XL U1048 ( .B0(n1925), .B1(n2246), .A0N(\register[25][29] ), .A1N(
        n2248), .Y(n303) );
  OAI2BB2XL U1049 ( .B0(n1922), .B1(n2246), .A0N(\register[25][30] ), .A1N(
        n2248), .Y(n304) );
  OAI2BB2XL U1050 ( .B0(n1919), .B1(n2246), .A0N(\register[25][31] ), .A1N(
        n2248), .Y(n305) );
  OAI2BB2XL U1051 ( .B0(n2012), .B1(n2242), .A0N(\register[24][0] ), .A1N(
        n2244), .Y(n306) );
  OAI2BB2XL U1052 ( .B0(n2009), .B1(n2242), .A0N(\register[24][1] ), .A1N(
        n2245), .Y(n307) );
  OAI2BB2XL U1053 ( .B0(n2006), .B1(n2242), .A0N(\register[24][2] ), .A1N(
        n2245), .Y(n308) );
  OAI2BB2XL U1054 ( .B0(n2003), .B1(n2242), .A0N(\register[24][3] ), .A1N(
        n2245), .Y(n309) );
  OAI2BB2XL U1055 ( .B0(n2000), .B1(n2242), .A0N(\register[24][4] ), .A1N(
        n2245), .Y(n310) );
  OAI2BB2XL U1056 ( .B0(n1997), .B1(n2242), .A0N(\register[24][5] ), .A1N(
        n2245), .Y(n311) );
  OAI2BB2XL U1057 ( .B0(n1994), .B1(n2242), .A0N(\register[24][6] ), .A1N(
        n2245), .Y(n312) );
  OAI2BB2XL U1058 ( .B0(n1991), .B1(n2242), .A0N(\register[24][7] ), .A1N(
        n2245), .Y(n313) );
  OAI2BB2XL U1059 ( .B0(n1988), .B1(n2243), .A0N(\register[24][8] ), .A1N(
        n2245), .Y(n314) );
  OAI2BB2XL U1060 ( .B0(n1985), .B1(n2243), .A0N(\register[24][9] ), .A1N(
        n2245), .Y(n315) );
  OAI2BB2XL U1061 ( .B0(n1982), .B1(n2243), .A0N(\register[24][10] ), .A1N(
        n2245), .Y(n316) );
  OAI2BB2XL U1062 ( .B0(n1979), .B1(n2243), .A0N(\register[24][11] ), .A1N(
        n2245), .Y(n317) );
  OAI2BB2XL U1063 ( .B0(n1976), .B1(n2243), .A0N(\register[24][12] ), .A1N(
        n2245), .Y(n318) );
  OAI2BB2XL U1064 ( .B0(n1973), .B1(n2243), .A0N(\register[24][13] ), .A1N(
        n2245), .Y(n319) );
  OAI2BB2XL U1065 ( .B0(n1970), .B1(n2243), .A0N(\register[24][14] ), .A1N(
        n2245), .Y(n320) );
  OAI2BB2XL U1066 ( .B0(n1967), .B1(n2243), .A0N(\register[24][15] ), .A1N(
        n2245), .Y(n321) );
  OAI2BB2XL U1067 ( .B0(n1964), .B1(n2244), .A0N(\register[24][16] ), .A1N(
        n2245), .Y(n322) );
  OAI2BB2XL U1068 ( .B0(n1961), .B1(n2244), .A0N(\register[24][17] ), .A1N(
        n2245), .Y(n323) );
  OAI2BB2XL U1069 ( .B0(n1958), .B1(n2243), .A0N(\register[24][18] ), .A1N(
        n2245), .Y(n324) );
  OAI2BB2XL U1070 ( .B0(n1955), .B1(n2244), .A0N(\register[24][19] ), .A1N(
        n2245), .Y(n325) );
  OAI2BB2XL U1071 ( .B0(n1952), .B1(n2244), .A0N(\register[24][20] ), .A1N(
        n2245), .Y(n326) );
  OAI2BB2XL U1072 ( .B0(n1949), .B1(n2244), .A0N(\register[24][21] ), .A1N(
        n2244), .Y(n327) );
  OAI2BB2XL U1073 ( .B0(n1946), .B1(n2244), .A0N(\register[24][22] ), .A1N(
        n2244), .Y(n328) );
  OAI2BB2XL U1074 ( .B0(n1943), .B1(n2244), .A0N(\register[24][23] ), .A1N(
        n2244), .Y(n329) );
  OAI2BB2XL U1075 ( .B0(n1940), .B1(n2244), .A0N(\register[24][24] ), .A1N(
        n2244), .Y(n330) );
  OAI2BB2XL U1076 ( .B0(n1937), .B1(n2243), .A0N(\register[24][25] ), .A1N(
        n2244), .Y(n331) );
  OAI2BB2XL U1077 ( .B0(n1934), .B1(n2243), .A0N(\register[24][26] ), .A1N(
        n2244), .Y(n332) );
  OAI2BB2XL U1078 ( .B0(n1931), .B1(n2243), .A0N(\register[24][27] ), .A1N(
        n2244), .Y(n333) );
  OAI2BB2XL U1079 ( .B0(n1928), .B1(n2242), .A0N(\register[24][28] ), .A1N(
        n2244), .Y(n334) );
  OAI2BB2XL U1080 ( .B0(n1925), .B1(n2242), .A0N(\register[24][29] ), .A1N(
        n2244), .Y(n335) );
  OAI2BB2XL U1081 ( .B0(n1922), .B1(n2242), .A0N(\register[24][30] ), .A1N(
        n2244), .Y(n336) );
  OAI2BB2XL U1082 ( .B0(n1919), .B1(n2242), .A0N(\register[24][31] ), .A1N(
        n2244), .Y(n337) );
  OAI2BB2XL U1083 ( .B0(n2011), .B1(n2206), .A0N(\register[15][0] ), .A1N(
        n2208), .Y(n594) );
  OAI2BB2XL U1084 ( .B0(n2008), .B1(n2206), .A0N(\register[15][1] ), .A1N(
        n2209), .Y(n595) );
  OAI2BB2XL U1085 ( .B0(n2005), .B1(n2206), .A0N(\register[15][2] ), .A1N(
        n2209), .Y(n596) );
  OAI2BB2XL U1086 ( .B0(n1963), .B1(n2208), .A0N(\register[15][16] ), .A1N(
        n2209), .Y(n610) );
  OAI2BB2XL U1087 ( .B0(n1960), .B1(n2208), .A0N(\register[15][17] ), .A1N(
        n2209), .Y(n611) );
  OAI2BB2XL U1088 ( .B0(n1957), .B1(n2207), .A0N(\register[15][18] ), .A1N(
        n2209), .Y(n612) );
  OAI2BB2XL U1089 ( .B0(n1954), .B1(n2208), .A0N(\register[15][19] ), .A1N(
        n2209), .Y(n613) );
  OAI2BB2XL U1090 ( .B0(n1951), .B1(n2208), .A0N(\register[15][20] ), .A1N(
        n2209), .Y(n614) );
  OAI2BB2XL U1091 ( .B0(n1948), .B1(n2208), .A0N(\register[15][21] ), .A1N(
        n2208), .Y(n615) );
  OAI2BB2XL U1092 ( .B0(n1945), .B1(n2208), .A0N(\register[15][22] ), .A1N(
        n2208), .Y(n616) );
  OAI2BB2XL U1093 ( .B0(n1942), .B1(n2208), .A0N(\register[15][23] ), .A1N(
        n2208), .Y(n617) );
  OAI2BB2XL U1094 ( .B0(n1939), .B1(n2208), .A0N(\register[15][24] ), .A1N(
        n2208), .Y(n618) );
  OAI2BB2XL U1095 ( .B0(n1936), .B1(n2207), .A0N(\register[15][25] ), .A1N(
        n2208), .Y(n619) );
  OAI2BB2XL U1096 ( .B0(n1933), .B1(n2207), .A0N(\register[15][26] ), .A1N(
        n2208), .Y(n620) );
  OAI2BB2XL U1097 ( .B0(n1930), .B1(n2207), .A0N(\register[15][27] ), .A1N(
        n2208), .Y(n621) );
  OAI2BB2XL U1098 ( .B0(n1927), .B1(n2206), .A0N(\register[15][28] ), .A1N(
        n2208), .Y(n622) );
  OAI2BB2XL U1099 ( .B0(n1924), .B1(n2206), .A0N(\register[15][29] ), .A1N(
        n2208), .Y(n623) );
  OAI2BB2XL U1100 ( .B0(n1921), .B1(n2206), .A0N(\register[15][30] ), .A1N(
        n2208), .Y(n624) );
  OAI2BB2XL U1101 ( .B0(n1918), .B1(n2206), .A0N(\register[15][31] ), .A1N(
        n2208), .Y(n625) );
  OAI2BB2XL U1102 ( .B0(n2011), .B1(n2202), .A0N(\register[14][0] ), .A1N(
        n2204), .Y(n626) );
  OAI2BB2XL U1103 ( .B0(n2008), .B1(n2202), .A0N(\register[14][1] ), .A1N(
        n2205), .Y(n627) );
  OAI2BB2XL U1104 ( .B0(n2002), .B1(n2202), .A0N(\register[14][3] ), .A1N(
        n2205), .Y(n629) );
  OAI2BB2XL U1105 ( .B0(n1999), .B1(n2202), .A0N(\register[14][4] ), .A1N(
        n2205), .Y(n630) );
  OAI2BB2XL U1106 ( .B0(n1996), .B1(n2202), .A0N(\register[14][5] ), .A1N(
        n2205), .Y(n631) );
  OAI2BB2XL U1107 ( .B0(n1993), .B1(n2202), .A0N(\register[14][6] ), .A1N(
        n2205), .Y(n632) );
  OAI2BB2XL U1108 ( .B0(n1990), .B1(n2202), .A0N(\register[14][7] ), .A1N(
        n2205), .Y(n633) );
  OAI2BB2XL U1109 ( .B0(n1987), .B1(n2203), .A0N(\register[14][8] ), .A1N(
        n2205), .Y(n634) );
  OAI2BB2XL U1110 ( .B0(n1984), .B1(n2203), .A0N(\register[14][9] ), .A1N(
        n2205), .Y(n635) );
  OAI2BB2XL U1111 ( .B0(n1981), .B1(n2203), .A0N(\register[14][10] ), .A1N(
        n2205), .Y(n636) );
  OAI2BB2XL U1112 ( .B0(n1978), .B1(n2203), .A0N(\register[14][11] ), .A1N(
        n2205), .Y(n637) );
  OAI2BB2XL U1113 ( .B0(n1975), .B1(n2203), .A0N(\register[14][12] ), .A1N(
        n2205), .Y(n638) );
  OAI2BB2XL U1114 ( .B0(n1972), .B1(n2203), .A0N(\register[14][13] ), .A1N(
        n2205), .Y(n639) );
  OAI2BB2XL U1115 ( .B0(n1969), .B1(n2203), .A0N(\register[14][14] ), .A1N(
        n2205), .Y(n640) );
  OAI2BB2XL U1116 ( .B0(n1966), .B1(n2203), .A0N(\register[14][15] ), .A1N(
        n2205), .Y(n641) );
  OAI2BB2XL U1117 ( .B0(n1963), .B1(n2204), .A0N(\register[14][16] ), .A1N(
        n2205), .Y(n642) );
  OAI2BB2XL U1118 ( .B0(n1960), .B1(n2204), .A0N(\register[14][17] ), .A1N(
        n2205), .Y(n643) );
  OAI2BB2XL U1119 ( .B0(n1957), .B1(n2203), .A0N(\register[14][18] ), .A1N(
        n2205), .Y(n644) );
  OAI2BB2XL U1120 ( .B0(n1954), .B1(n2204), .A0N(\register[14][19] ), .A1N(
        n2205), .Y(n645) );
  OAI2BB2XL U1121 ( .B0(n1951), .B1(n2204), .A0N(\register[14][20] ), .A1N(
        n2205), .Y(n646) );
  OAI2BB2XL U1122 ( .B0(n1948), .B1(n2204), .A0N(\register[14][21] ), .A1N(
        n2204), .Y(n647) );
  OAI2BB2XL U1123 ( .B0(n1945), .B1(n2204), .A0N(\register[14][22] ), .A1N(
        n2204), .Y(n648) );
  OAI2BB2XL U1124 ( .B0(n1942), .B1(n2204), .A0N(\register[14][23] ), .A1N(
        n2204), .Y(n649) );
  OAI2BB2XL U1125 ( .B0(n1939), .B1(n2204), .A0N(\register[14][24] ), .A1N(
        n2204), .Y(n650) );
  OAI2BB2XL U1126 ( .B0(n1936), .B1(n2203), .A0N(\register[14][25] ), .A1N(
        n2204), .Y(n651) );
  OAI2BB2XL U1127 ( .B0(n1933), .B1(n2203), .A0N(\register[14][26] ), .A1N(
        n2204), .Y(n652) );
  OAI2BB2XL U1128 ( .B0(n1930), .B1(n2203), .A0N(\register[14][27] ), .A1N(
        n2204), .Y(n653) );
  OAI2BB2XL U1129 ( .B0(n1927), .B1(n2202), .A0N(\register[14][28] ), .A1N(
        n2204), .Y(n654) );
  OAI2BB2XL U1130 ( .B0(n1924), .B1(n2202), .A0N(\register[14][29] ), .A1N(
        n2204), .Y(n655) );
  OAI2BB2XL U1131 ( .B0(n1921), .B1(n2202), .A0N(\register[14][30] ), .A1N(
        n2204), .Y(n656) );
  OAI2BB2XL U1132 ( .B0(n1918), .B1(n2202), .A0N(\register[14][31] ), .A1N(
        n2204), .Y(n657) );
  OAI2BB2XL U1133 ( .B0(n2011), .B1(n2198), .A0N(\register[13][0] ), .A1N(
        n2200), .Y(n658) );
  OAI2BB2XL U1134 ( .B0(n2008), .B1(n2198), .A0N(\register[13][1] ), .A1N(
        n2201), .Y(n659) );
  OAI2BB2XL U1135 ( .B0(n2005), .B1(n2198), .A0N(\register[13][2] ), .A1N(
        n2201), .Y(n660) );
  OAI2BB2XL U1136 ( .B0(n2002), .B1(n2198), .A0N(\register[13][3] ), .A1N(
        n2201), .Y(n661) );
  OAI2BB2XL U1137 ( .B0(n1999), .B1(n2198), .A0N(\register[13][4] ), .A1N(
        n2201), .Y(n662) );
  OAI2BB2XL U1138 ( .B0(n1996), .B1(n2198), .A0N(\register[13][5] ), .A1N(
        n2201), .Y(n663) );
  OAI2BB2XL U1139 ( .B0(n1993), .B1(n2198), .A0N(\register[13][6] ), .A1N(
        n2201), .Y(n664) );
  OAI2BB2XL U1140 ( .B0(n1990), .B1(n2198), .A0N(\register[13][7] ), .A1N(
        n2201), .Y(n665) );
  OAI2BB2XL U1141 ( .B0(n1987), .B1(n2199), .A0N(\register[13][8] ), .A1N(
        n2201), .Y(n666) );
  OAI2BB2XL U1142 ( .B0(n1981), .B1(n2199), .A0N(\register[13][10] ), .A1N(
        n2201), .Y(n668) );
  OAI2BB2XL U1143 ( .B0(n1978), .B1(n2199), .A0N(\register[13][11] ), .A1N(
        n2201), .Y(n669) );
  OAI2BB2XL U1144 ( .B0(n1975), .B1(n2199), .A0N(\register[13][12] ), .A1N(
        n2201), .Y(n670) );
  OAI2BB2XL U1145 ( .B0(n1972), .B1(n2199), .A0N(\register[13][13] ), .A1N(
        n2201), .Y(n671) );
  OAI2BB2XL U1146 ( .B0(n1969), .B1(n2199), .A0N(\register[13][14] ), .A1N(
        n2201), .Y(n672) );
  OAI2BB2XL U1147 ( .B0(n1966), .B1(n2199), .A0N(\register[13][15] ), .A1N(
        n2201), .Y(n673) );
  OAI2BB2XL U1148 ( .B0(n1963), .B1(n2200), .A0N(\register[13][16] ), .A1N(
        n2201), .Y(n674) );
  OAI2BB2XL U1149 ( .B0(n1960), .B1(n2200), .A0N(\register[13][17] ), .A1N(
        n2201), .Y(n675) );
  OAI2BB2XL U1150 ( .B0(n1957), .B1(n2199), .A0N(\register[13][18] ), .A1N(
        n2201), .Y(n676) );
  OAI2BB2XL U1151 ( .B0(n1954), .B1(n2200), .A0N(\register[13][19] ), .A1N(
        n2201), .Y(n677) );
  OAI2BB2XL U1152 ( .B0(n1951), .B1(n2200), .A0N(\register[13][20] ), .A1N(
        n2201), .Y(n678) );
  OAI2BB2XL U1153 ( .B0(n1948), .B1(n2200), .A0N(\register[13][21] ), .A1N(
        n2200), .Y(n679) );
  OAI2BB2XL U1154 ( .B0(n1945), .B1(n2200), .A0N(\register[13][22] ), .A1N(
        n2200), .Y(n680) );
  OAI2BB2XL U1155 ( .B0(n1942), .B1(n2200), .A0N(\register[13][23] ), .A1N(
        n2200), .Y(n681) );
  OAI2BB2XL U1156 ( .B0(n1939), .B1(n2200), .A0N(\register[13][24] ), .A1N(
        n2200), .Y(n682) );
  OAI2BB2XL U1157 ( .B0(n1936), .B1(n2199), .A0N(\register[13][25] ), .A1N(
        n2200), .Y(n683) );
  OAI2BB2XL U1158 ( .B0(n1933), .B1(n2199), .A0N(\register[13][26] ), .A1N(
        n2200), .Y(n684) );
  OAI2BB2XL U1159 ( .B0(n1930), .B1(n2199), .A0N(\register[13][27] ), .A1N(
        n2200), .Y(n685) );
  OAI2BB2XL U1160 ( .B0(n1927), .B1(n2198), .A0N(\register[13][28] ), .A1N(
        n2200), .Y(n686) );
  OAI2BB2XL U1161 ( .B0(n1924), .B1(n2198), .A0N(\register[13][29] ), .A1N(
        n2200), .Y(n687) );
  OAI2BB2XL U1162 ( .B0(n1921), .B1(n2198), .A0N(\register[13][30] ), .A1N(
        n2200), .Y(n688) );
  OAI2BB2XL U1163 ( .B0(n1918), .B1(n2198), .A0N(\register[13][31] ), .A1N(
        n2200), .Y(n689) );
  OAI2BB2XL U1164 ( .B0(n2011), .B1(n2194), .A0N(\register[12][0] ), .A1N(
        n2196), .Y(n690) );
  OAI2BB2XL U1165 ( .B0(n2008), .B1(n2194), .A0N(\register[12][1] ), .A1N(
        n2197), .Y(n691) );
  OAI2BB2XL U1166 ( .B0(n2005), .B1(n2194), .A0N(\register[12][2] ), .A1N(
        n2197), .Y(n692) );
  OAI2BB2XL U1167 ( .B0(n2002), .B1(n2194), .A0N(\register[12][3] ), .A1N(
        n2197), .Y(n693) );
  OAI2BB2XL U1168 ( .B0(n1999), .B1(n2194), .A0N(\register[12][4] ), .A1N(
        n2197), .Y(n694) );
  OAI2BB2XL U1169 ( .B0(n1996), .B1(n2194), .A0N(\register[12][5] ), .A1N(
        n2197), .Y(n695) );
  OAI2BB2XL U1170 ( .B0(n1993), .B1(n2194), .A0N(\register[12][6] ), .A1N(
        n2197), .Y(n696) );
  OAI2BB2XL U1171 ( .B0(n1990), .B1(n2194), .A0N(\register[12][7] ), .A1N(
        n2197), .Y(n697) );
  OAI2BB2XL U1172 ( .B0(n1987), .B1(n2195), .A0N(\register[12][8] ), .A1N(
        n2197), .Y(n698) );
  OAI2BB2XL U1173 ( .B0(n1984), .B1(n2195), .A0N(\register[12][9] ), .A1N(
        n2197), .Y(n699) );
  OAI2BB2XL U1174 ( .B0(n1981), .B1(n2195), .A0N(\register[12][10] ), .A1N(
        n2197), .Y(n700) );
  OAI2BB2XL U1175 ( .B0(n1978), .B1(n2195), .A0N(\register[12][11] ), .A1N(
        n2197), .Y(n701) );
  OAI2BB2XL U1176 ( .B0(n1975), .B1(n2195), .A0N(\register[12][12] ), .A1N(
        n2197), .Y(n702) );
  OAI2BB2XL U1177 ( .B0(n1972), .B1(n2195), .A0N(\register[12][13] ), .A1N(
        n2197), .Y(n703) );
  OAI2BB2XL U1178 ( .B0(n1969), .B1(n2195), .A0N(\register[12][14] ), .A1N(
        n2197), .Y(n704) );
  OAI2BB2XL U1179 ( .B0(n1966), .B1(n2195), .A0N(\register[12][15] ), .A1N(
        n2197), .Y(n705) );
  OAI2BB2XL U1180 ( .B0(n1963), .B1(n2196), .A0N(\register[12][16] ), .A1N(
        n2197), .Y(n706) );
  OAI2BB2XL U1181 ( .B0(n1960), .B1(n2196), .A0N(\register[12][17] ), .A1N(
        n2197), .Y(n707) );
  OAI2BB2XL U1182 ( .B0(n1957), .B1(n2195), .A0N(\register[12][18] ), .A1N(
        n2197), .Y(n708) );
  OAI2BB2XL U1183 ( .B0(n1954), .B1(n2196), .A0N(\register[12][19] ), .A1N(
        n2197), .Y(n709) );
  OAI2BB2XL U1184 ( .B0(n1951), .B1(n2196), .A0N(\register[12][20] ), .A1N(
        n2197), .Y(n710) );
  OAI2BB2XL U1185 ( .B0(n1948), .B1(n2196), .A0N(\register[12][21] ), .A1N(
        n2196), .Y(n711) );
  OAI2BB2XL U1186 ( .B0(n1945), .B1(n2196), .A0N(\register[12][22] ), .A1N(
        n2196), .Y(n712) );
  OAI2BB2XL U1187 ( .B0(n1942), .B1(n2196), .A0N(\register[12][23] ), .A1N(
        n2196), .Y(n713) );
  OAI2BB2XL U1188 ( .B0(n1939), .B1(n2196), .A0N(\register[12][24] ), .A1N(
        n2196), .Y(n714) );
  OAI2BB2XL U1189 ( .B0(n1936), .B1(n2195), .A0N(\register[12][25] ), .A1N(
        n2196), .Y(n715) );
  OAI2BB2XL U1190 ( .B0(n1933), .B1(n2195), .A0N(\register[12][26] ), .A1N(
        n2196), .Y(n716) );
  OAI2BB2XL U1191 ( .B0(n1930), .B1(n2195), .A0N(\register[12][27] ), .A1N(
        n2196), .Y(n717) );
  OAI2BB2XL U1192 ( .B0(n1927), .B1(n2194), .A0N(\register[12][28] ), .A1N(
        n2196), .Y(n718) );
  OAI2BB2XL U1193 ( .B0(n1924), .B1(n2194), .A0N(\register[12][29] ), .A1N(
        n2196), .Y(n719) );
  OAI2BB2XL U1194 ( .B0(n1921), .B1(n2194), .A0N(\register[12][30] ), .A1N(
        n2196), .Y(n720) );
  OAI2BB2XL U1195 ( .B0(n1918), .B1(n2194), .A0N(\register[12][31] ), .A1N(
        n2196), .Y(n721) );
  OAI2BB2XL U1196 ( .B0(n2010), .B1(n2190), .A0N(\register[11][0] ), .A1N(
        n2192), .Y(n722) );
  OAI2BB2XL U1197 ( .B0(n2007), .B1(n2190), .A0N(\register[11][1] ), .A1N(
        n2193), .Y(n723) );
  OAI2BB2XL U1198 ( .B0(n2004), .B1(n2190), .A0N(\register[11][2] ), .A1N(
        n2193), .Y(n724) );
  OAI2BB2XL U1199 ( .B0(n2001), .B1(n2190), .A0N(\register[11][3] ), .A1N(
        n2193), .Y(n725) );
  OAI2BB2XL U1200 ( .B0(n1998), .B1(n2190), .A0N(\register[11][4] ), .A1N(
        n2193), .Y(n726) );
  OAI2BB2XL U1201 ( .B0(n1995), .B1(n2190), .A0N(\register[11][5] ), .A1N(
        n2193), .Y(n727) );
  OAI2BB2XL U1202 ( .B0(n1983), .B1(n2191), .A0N(\register[11][9] ), .A1N(
        n2193), .Y(n731) );
  OAI2BB2XL U1203 ( .B0(n1980), .B1(n2191), .A0N(\register[11][10] ), .A1N(
        n2193), .Y(n732) );
  OAI2BB2XL U1204 ( .B0(n1977), .B1(n2191), .A0N(\register[11][11] ), .A1N(
        n2193), .Y(n733) );
  OAI2BB2XL U1205 ( .B0(n1974), .B1(n2191), .A0N(\register[11][12] ), .A1N(
        n2193), .Y(n734) );
  OAI2BB2XL U1206 ( .B0(n1971), .B1(n2191), .A0N(\register[11][13] ), .A1N(
        n2193), .Y(n735) );
  OAI2BB2XL U1207 ( .B0(n1968), .B1(n2191), .A0N(\register[11][14] ), .A1N(
        n2193), .Y(n736) );
  OAI2BB2XL U1208 ( .B0(n1965), .B1(n2191), .A0N(\register[11][15] ), .A1N(
        n2193), .Y(n737) );
  OAI2BB2XL U1209 ( .B0(n1962), .B1(n2192), .A0N(\register[11][16] ), .A1N(
        n2193), .Y(n738) );
  OAI2BB2XL U1210 ( .B0(n1959), .B1(n2192), .A0N(\register[11][17] ), .A1N(
        n2193), .Y(n739) );
  OAI2BB2XL U1211 ( .B0(n1956), .B1(n2191), .A0N(\register[11][18] ), .A1N(
        n2193), .Y(n740) );
  OAI2BB2XL U1212 ( .B0(n1953), .B1(n2192), .A0N(\register[11][19] ), .A1N(
        n2193), .Y(n741) );
  OAI2BB2XL U1213 ( .B0(n1950), .B1(n2192), .A0N(\register[11][20] ), .A1N(
        n2193), .Y(n742) );
  OAI2BB2XL U1214 ( .B0(n1947), .B1(n2192), .A0N(\register[11][21] ), .A1N(
        n2192), .Y(n743) );
  OAI2BB2XL U1215 ( .B0(n1944), .B1(n2192), .A0N(\register[11][22] ), .A1N(
        n2192), .Y(n744) );
  OAI2BB2XL U1216 ( .B0(n1941), .B1(n2192), .A0N(\register[11][23] ), .A1N(
        n2192), .Y(n745) );
  OAI2BB2XL U1217 ( .B0(n1938), .B1(n2192), .A0N(\register[11][24] ), .A1N(
        n2192), .Y(n746) );
  OAI2BB2XL U1218 ( .B0(n1935), .B1(n2191), .A0N(\register[11][25] ), .A1N(
        n2192), .Y(n747) );
  OAI2BB2XL U1219 ( .B0(n1932), .B1(n2191), .A0N(\register[11][26] ), .A1N(
        n2192), .Y(n748) );
  OAI2BB2XL U1220 ( .B0(n1929), .B1(n2191), .A0N(\register[11][27] ), .A1N(
        n2192), .Y(n749) );
  OAI2BB2XL U1221 ( .B0(n1926), .B1(n2190), .A0N(\register[11][28] ), .A1N(
        n2192), .Y(n750) );
  OAI2BB2XL U1222 ( .B0(n1923), .B1(n2190), .A0N(\register[11][29] ), .A1N(
        n2192), .Y(n751) );
  OAI2BB2XL U1223 ( .B0(n1920), .B1(n2190), .A0N(\register[11][30] ), .A1N(
        n2192), .Y(n752) );
  OAI2BB2XL U1224 ( .B0(n1950), .B1(n2188), .A0N(\register[10][20] ), .A1N(
        n2189), .Y(n774) );
  OAI2BB2XL U1225 ( .B0(n1947), .B1(n2188), .A0N(\register[10][21] ), .A1N(
        n2188), .Y(n775) );
  OAI2BB2XL U1226 ( .B0(n1944), .B1(n2188), .A0N(\register[10][22] ), .A1N(
        n2188), .Y(n776) );
  OAI2BB2XL U1227 ( .B0(n1941), .B1(n2188), .A0N(\register[10][23] ), .A1N(
        n2188), .Y(n777) );
  OAI2BB2XL U1228 ( .B0(n1938), .B1(n2188), .A0N(\register[10][24] ), .A1N(
        n2188), .Y(n778) );
  OAI2BB2XL U1229 ( .B0(n2010), .B1(n2182), .A0N(\register[9][0] ), .A1N(n2184), .Y(n786) );
  OAI2BB2XL U1230 ( .B0(n2007), .B1(n2182), .A0N(\register[9][1] ), .A1N(n2185), .Y(n787) );
  OAI2BB2XL U1231 ( .B0(n1998), .B1(n2182), .A0N(\register[9][4] ), .A1N(n2185), .Y(n790) );
  OAI2BB2XL U1232 ( .B0(n1995), .B1(n2182), .A0N(\register[9][5] ), .A1N(n2185), .Y(n791) );
  OAI2BB2XL U1233 ( .B0(n1992), .B1(n2182), .A0N(\register[9][6] ), .A1N(n2185), .Y(n792) );
  OAI2BB2XL U1234 ( .B0(n1989), .B1(n2182), .A0N(\register[9][7] ), .A1N(n2185), .Y(n793) );
  OAI2BB2XL U1235 ( .B0(n1986), .B1(n2183), .A0N(\register[9][8] ), .A1N(n2185), .Y(n794) );
  OAI2BB2XL U1236 ( .B0(n1983), .B1(n2183), .A0N(\register[9][9] ), .A1N(n2185), .Y(n795) );
  OAI2BB2XL U1237 ( .B0(n1980), .B1(n2183), .A0N(\register[9][10] ), .A1N(
        n2185), .Y(n796) );
  OAI2BB2XL U1238 ( .B0(n1977), .B1(n2183), .A0N(\register[9][11] ), .A1N(
        n2185), .Y(n797) );
  OAI2BB2XL U1239 ( .B0(n1974), .B1(n2183), .A0N(\register[9][12] ), .A1N(
        n2185), .Y(n798) );
  OAI2BB2XL U1240 ( .B0(n1971), .B1(n2183), .A0N(\register[9][13] ), .A1N(
        n2185), .Y(n799) );
  OAI2BB2XL U1241 ( .B0(n1968), .B1(n2183), .A0N(\register[9][14] ), .A1N(
        n2185), .Y(n800) );
  OAI2BB2XL U1242 ( .B0(n1965), .B1(n2183), .A0N(\register[9][15] ), .A1N(
        n2185), .Y(n801) );
  OAI2BB2XL U1243 ( .B0(n1959), .B1(n2184), .A0N(\register[9][17] ), .A1N(
        n2185), .Y(n803) );
  OAI2BB2XL U1244 ( .B0(n1953), .B1(n2184), .A0N(\register[9][19] ), .A1N(
        n2185), .Y(n805) );
  OAI2BB2XL U1245 ( .B0(n1950), .B1(n2184), .A0N(\register[9][20] ), .A1N(
        n2185), .Y(n806) );
  OAI2BB2XL U1246 ( .B0(n1947), .B1(n2184), .A0N(\register[9][21] ), .A1N(
        n2184), .Y(n807) );
  OAI2BB2XL U1247 ( .B0(n1944), .B1(n2184), .A0N(\register[9][22] ), .A1N(
        n2184), .Y(n808) );
  OAI2BB2XL U1248 ( .B0(n1941), .B1(n2184), .A0N(\register[9][23] ), .A1N(
        n2184), .Y(n809) );
  OAI2BB2XL U1249 ( .B0(n1938), .B1(n2184), .A0N(\register[9][24] ), .A1N(
        n2184), .Y(n810) );
  OAI2BB2XL U1250 ( .B0(n2010), .B1(n2178), .A0N(\register[8][0] ), .A1N(n2180), .Y(n818) );
  OAI2BB2XL U1251 ( .B0(n2007), .B1(n2178), .A0N(\register[8][1] ), .A1N(n2181), .Y(n819) );
  OAI2BB2XL U1252 ( .B0(n2004), .B1(n2178), .A0N(\register[8][2] ), .A1N(n2181), .Y(n820) );
  OAI2BB2XL U1253 ( .B0(n2001), .B1(n2178), .A0N(\register[8][3] ), .A1N(n2181), .Y(n821) );
  OAI2BB2XL U1254 ( .B0(n1998), .B1(n2178), .A0N(\register[8][4] ), .A1N(n2181), .Y(n822) );
  OAI2BB2XL U1255 ( .B0(n1995), .B1(n2178), .A0N(\register[8][5] ), .A1N(n2181), .Y(n823) );
  OAI2BB2XL U1256 ( .B0(n1992), .B1(n2178), .A0N(\register[8][6] ), .A1N(n2181), .Y(n824) );
  OAI2BB2XL U1257 ( .B0(n1989), .B1(n2178), .A0N(\register[8][7] ), .A1N(n2181), .Y(n825) );
  OAI2BB2XL U1258 ( .B0(n1986), .B1(n2179), .A0N(\register[8][8] ), .A1N(n2181), .Y(n826) );
  OAI2BB2XL U1259 ( .B0(n1983), .B1(n2179), .A0N(\register[8][9] ), .A1N(n2181), .Y(n827) );
  OAI2BB2XL U1260 ( .B0(n1980), .B1(n2179), .A0N(\register[8][10] ), .A1N(
        n2181), .Y(n828) );
  OAI2BB2XL U1261 ( .B0(n1977), .B1(n2179), .A0N(\register[8][11] ), .A1N(
        n2181), .Y(n829) );
  OAI2BB2XL U1262 ( .B0(n1974), .B1(n2179), .A0N(\register[8][12] ), .A1N(
        n2181), .Y(n830) );
  OAI2BB2XL U1263 ( .B0(n1971), .B1(n2179), .A0N(\register[8][13] ), .A1N(
        n2181), .Y(n831) );
  OAI2BB2XL U1264 ( .B0(n1968), .B1(n2179), .A0N(\register[8][14] ), .A1N(
        n2181), .Y(n832) );
  OAI2BB2XL U1265 ( .B0(n1965), .B1(n2179), .A0N(\register[8][15] ), .A1N(
        n2181), .Y(n833) );
  OAI2BB2XL U1266 ( .B0(n1962), .B1(n2180), .A0N(\register[8][16] ), .A1N(
        n2181), .Y(n834) );
  OAI2BB2XL U1267 ( .B0(n1959), .B1(n2180), .A0N(\register[8][17] ), .A1N(
        n2181), .Y(n835) );
  OAI2BB2XL U1268 ( .B0(n1956), .B1(n2179), .A0N(\register[8][18] ), .A1N(
        n2181), .Y(n836) );
  OAI2BB2XL U1269 ( .B0(n1953), .B1(n2180), .A0N(\register[8][19] ), .A1N(
        n2181), .Y(n837) );
  OAI2BB2XL U1270 ( .B0(n1950), .B1(n2180), .A0N(\register[8][20] ), .A1N(
        n2181), .Y(n838) );
  OAI2BB2XL U1271 ( .B0(n1947), .B1(n2180), .A0N(\register[8][21] ), .A1N(
        n2180), .Y(n839) );
  OAI2BB2XL U1272 ( .B0(n1944), .B1(n2180), .A0N(\register[8][22] ), .A1N(
        n2180), .Y(n840) );
  OAI2BB2XL U1273 ( .B0(n1941), .B1(n2180), .A0N(\register[8][23] ), .A1N(
        n2180), .Y(n841) );
  OAI2BB2XL U1274 ( .B0(n1938), .B1(n2180), .A0N(\register[8][24] ), .A1N(
        n2180), .Y(n842) );
  OAI2BB2XL U1275 ( .B0(n1923), .B1(n2178), .A0N(\register[8][29] ), .A1N(
        n2180), .Y(n847) );
  OAI2BB2XL U1276 ( .B0(n1917), .B1(n2178), .A0N(\register[8][31] ), .A1N(
        n2180), .Y(n849) );
  OAI2BB2XL U1277 ( .B0(n2010), .B1(n2174), .A0N(\register[7][0] ), .A1N(n2176), .Y(n850) );
  OAI2BB2XL U1278 ( .B0(n2007), .B1(n2174), .A0N(\register[7][1] ), .A1N(n2177), .Y(n851) );
  OAI2BB2XL U1279 ( .B0(n2004), .B1(n2174), .A0N(\register[7][2] ), .A1N(n2177), .Y(n852) );
  OAI2BB2XL U1280 ( .B0(n2001), .B1(n2174), .A0N(\register[7][3] ), .A1N(n2177), .Y(n853) );
  OAI2BB2XL U1281 ( .B0(n1998), .B1(n2174), .A0N(\register[7][4] ), .A1N(n2177), .Y(n854) );
  OAI2BB2XL U1282 ( .B0(n1995), .B1(n2174), .A0N(\register[7][5] ), .A1N(n2177), .Y(n855) );
  OAI2BB2XL U1283 ( .B0(n1992), .B1(n2174), .A0N(\register[7][6] ), .A1N(n2177), .Y(n856) );
  OAI2BB2XL U1284 ( .B0(n1989), .B1(n2174), .A0N(\register[7][7] ), .A1N(n2177), .Y(n857) );
  OAI2BB2XL U1285 ( .B0(n1986), .B1(n2175), .A0N(\register[7][8] ), .A1N(n2177), .Y(n858) );
  OAI2BB2XL U1286 ( .B0(n1983), .B1(n2175), .A0N(\register[7][9] ), .A1N(n2177), .Y(n859) );
  OAI2BB2XL U1287 ( .B0(n1980), .B1(n2175), .A0N(\register[7][10] ), .A1N(
        n2177), .Y(n860) );
  OAI2BB2XL U1288 ( .B0(n1977), .B1(n2175), .A0N(\register[7][11] ), .A1N(
        n2177), .Y(n861) );
  OAI2BB2XL U1289 ( .B0(n1974), .B1(n2175), .A0N(\register[7][12] ), .A1N(
        n2177), .Y(n862) );
  OAI2BB2XL U1290 ( .B0(n1971), .B1(n2175), .A0N(\register[7][13] ), .A1N(
        n2177), .Y(n863) );
  OAI2BB2XL U1291 ( .B0(n1965), .B1(n2175), .A0N(\register[7][15] ), .A1N(
        n2177), .Y(n865) );
  OAI2BB2XL U1292 ( .B0(n1962), .B1(n2176), .A0N(\register[7][16] ), .A1N(
        n2177), .Y(n866) );
  OAI2BB2XL U1293 ( .B0(n1953), .B1(n2176), .A0N(\register[7][19] ), .A1N(
        n2177), .Y(n869) );
  OAI2BB2XL U1294 ( .B0(n1950), .B1(n2176), .A0N(\register[7][20] ), .A1N(
        n2177), .Y(n870) );
  OAI2BB2XL U1295 ( .B0(n1947), .B1(n2176), .A0N(\register[7][21] ), .A1N(
        n2176), .Y(n871) );
  OAI2BB2XL U1296 ( .B0(n1929), .B1(n2175), .A0N(\register[7][27] ), .A1N(
        n2176), .Y(n877) );
  OAI2BB2XL U1297 ( .B0(n1926), .B1(n2174), .A0N(\register[7][28] ), .A1N(
        n2176), .Y(n878) );
  OAI2BB2XL U1298 ( .B0(n1923), .B1(n2174), .A0N(\register[7][29] ), .A1N(
        n2176), .Y(n879) );
  OAI2BB2XL U1299 ( .B0(n1920), .B1(n2174), .A0N(\register[7][30] ), .A1N(
        n2176), .Y(n880) );
  OAI2BB2XL U1300 ( .B0(n1917), .B1(n2174), .A0N(\register[7][31] ), .A1N(
        n2176), .Y(n881) );
  OAI2BB2XL U1301 ( .B0(n2010), .B1(n2170), .A0N(\register[6][0] ), .A1N(n2172), .Y(n882) );
  OAI2BB2XL U1302 ( .B0(n2007), .B1(n2170), .A0N(\register[6][1] ), .A1N(n2173), .Y(n883) );
  OAI2BB2XL U1303 ( .B0(n2004), .B1(n2170), .A0N(\register[6][2] ), .A1N(n2173), .Y(n884) );
  OAI2BB2XL U1304 ( .B0(n2001), .B1(n2170), .A0N(\register[6][3] ), .A1N(n2173), .Y(n885) );
  OAI2BB2XL U1305 ( .B0(n1998), .B1(n2170), .A0N(\register[6][4] ), .A1N(n2173), .Y(n886) );
  OAI2BB2XL U1306 ( .B0(n1995), .B1(n2170), .A0N(\register[6][5] ), .A1N(n2173), .Y(n887) );
  OAI2BB2XL U1307 ( .B0(n1992), .B1(n2170), .A0N(\register[6][6] ), .A1N(n2173), .Y(n888) );
  OAI2BB2XL U1308 ( .B0(n1989), .B1(n2170), .A0N(\register[6][7] ), .A1N(n2173), .Y(n889) );
  OAI2BB2XL U1309 ( .B0(n1986), .B1(n2171), .A0N(\register[6][8] ), .A1N(n2173), .Y(n890) );
  OAI2BB2XL U1310 ( .B0(n1983), .B1(n2171), .A0N(\register[6][9] ), .A1N(n2173), .Y(n891) );
  OAI2BB2XL U1311 ( .B0(n1980), .B1(n2171), .A0N(\register[6][10] ), .A1N(
        n2173), .Y(n892) );
  OAI2BB2XL U1312 ( .B0(n1977), .B1(n2171), .A0N(\register[6][11] ), .A1N(
        n2173), .Y(n893) );
  OAI2BB2XL U1313 ( .B0(n1974), .B1(n2171), .A0N(\register[6][12] ), .A1N(
        n2173), .Y(n894) );
  OAI2BB2XL U1314 ( .B0(n1971), .B1(n2171), .A0N(\register[6][13] ), .A1N(
        n2173), .Y(n895) );
  OAI2BB2XL U1315 ( .B0(n1968), .B1(n2171), .A0N(\register[6][14] ), .A1N(
        n2173), .Y(n896) );
  OAI2BB2XL U1316 ( .B0(n1965), .B1(n2171), .A0N(\register[6][15] ), .A1N(
        n2173), .Y(n897) );
  OAI2BB2XL U1317 ( .B0(n1962), .B1(n2172), .A0N(\register[6][16] ), .A1N(
        n2173), .Y(n898) );
  OAI2BB2XL U1318 ( .B0(n1959), .B1(n2172), .A0N(\register[6][17] ), .A1N(
        n2173), .Y(n899) );
  OAI2BB2XL U1319 ( .B0(n1956), .B1(n2171), .A0N(\register[6][18] ), .A1N(
        n2173), .Y(n900) );
  OAI2BB2XL U1320 ( .B0(n1953), .B1(n2172), .A0N(\register[6][19] ), .A1N(
        n2173), .Y(n901) );
  OAI2BB2XL U1321 ( .B0(n1950), .B1(n2172), .A0N(\register[6][20] ), .A1N(
        n2173), .Y(n902) );
  OAI2BB2XL U1322 ( .B0(n1947), .B1(n2172), .A0N(\register[6][21] ), .A1N(
        n2172), .Y(n903) );
  OAI2BB2XL U1323 ( .B0(n1944), .B1(n2172), .A0N(\register[6][22] ), .A1N(
        n2172), .Y(n904) );
  OAI2BB2XL U1324 ( .B0(n1938), .B1(n2172), .A0N(\register[6][24] ), .A1N(
        n2172), .Y(n906) );
  OAI2BB2XL U1325 ( .B0(n1935), .B1(n2171), .A0N(\register[6][25] ), .A1N(
        n2172), .Y(n907) );
  OAI2BB2XL U1326 ( .B0(n1932), .B1(n2171), .A0N(\register[6][26] ), .A1N(
        n2172), .Y(n908) );
  OAI2BB2XL U1327 ( .B0(n1929), .B1(n2171), .A0N(\register[6][27] ), .A1N(
        n2172), .Y(n909) );
  OAI2BB2XL U1328 ( .B0(n1926), .B1(n2170), .A0N(\register[6][28] ), .A1N(
        n2172), .Y(n910) );
  OAI2BB2XL U1329 ( .B0(n1923), .B1(n2170), .A0N(\register[6][29] ), .A1N(
        n2172), .Y(n911) );
  OAI2BB2XL U1330 ( .B0(n1920), .B1(n2170), .A0N(\register[6][30] ), .A1N(
        n2172), .Y(n912) );
  OAI2BB2XL U1331 ( .B0(n1917), .B1(n2170), .A0N(\register[6][31] ), .A1N(
        n2172), .Y(n913) );
  OAI2BB2XL U1332 ( .B0(n2010), .B1(n2166), .A0N(\register[5][0] ), .A1N(n2168), .Y(n914) );
  OAI2BB2XL U1333 ( .B0(n2007), .B1(n2166), .A0N(\register[5][1] ), .A1N(n2169), .Y(n915) );
  OAI2BB2XL U1334 ( .B0(n2004), .B1(n2166), .A0N(\register[5][2] ), .A1N(n2169), .Y(n916) );
  OAI2BB2XL U1335 ( .B0(n2001), .B1(n2166), .A0N(\register[5][3] ), .A1N(n2169), .Y(n917) );
  OAI2BB2XL U1336 ( .B0(n1998), .B1(n2166), .A0N(\register[5][4] ), .A1N(n2169), .Y(n918) );
  OAI2BB2XL U1337 ( .B0(n1995), .B1(n2166), .A0N(\register[5][5] ), .A1N(n2169), .Y(n919) );
  OAI2BB2XL U1338 ( .B0(n1992), .B1(n2166), .A0N(\register[5][6] ), .A1N(n2169), .Y(n920) );
  OAI2BB2XL U1339 ( .B0(n1989), .B1(n2166), .A0N(\register[5][7] ), .A1N(n2169), .Y(n921) );
  OAI2BB2XL U1340 ( .B0(n1986), .B1(n2167), .A0N(\register[5][8] ), .A1N(n2169), .Y(n922) );
  OAI2BB2XL U1341 ( .B0(n1983), .B1(n2167), .A0N(\register[5][9] ), .A1N(n2169), .Y(n923) );
  OAI2BB2XL U1342 ( .B0(n1980), .B1(n2167), .A0N(\register[5][10] ), .A1N(
        n2169), .Y(n924) );
  OAI2BB2XL U1343 ( .B0(n1977), .B1(n2167), .A0N(\register[5][11] ), .A1N(
        n2169), .Y(n925) );
  OAI2BB2XL U1344 ( .B0(n1974), .B1(n2167), .A0N(\register[5][12] ), .A1N(
        n2169), .Y(n926) );
  OAI2BB2XL U1345 ( .B0(n1971), .B1(n2167), .A0N(\register[5][13] ), .A1N(
        n2169), .Y(n927) );
  OAI2BB2XL U1346 ( .B0(n1968), .B1(n2167), .A0N(\register[5][14] ), .A1N(
        n2169), .Y(n928) );
  OAI2BB2XL U1347 ( .B0(n1965), .B1(n2167), .A0N(\register[5][15] ), .A1N(
        n2169), .Y(n929) );
  OAI2BB2XL U1348 ( .B0(n1962), .B1(n2168), .A0N(\register[5][16] ), .A1N(
        n2169), .Y(n930) );
  OAI2BB2XL U1349 ( .B0(n1959), .B1(n2168), .A0N(\register[5][17] ), .A1N(
        n2169), .Y(n931) );
  OAI2BB2XL U1350 ( .B0(n1956), .B1(n2167), .A0N(\register[5][18] ), .A1N(
        n2169), .Y(n932) );
  OAI2BB2XL U1351 ( .B0(n1953), .B1(n2168), .A0N(\register[5][19] ), .A1N(
        n2169), .Y(n933) );
  OAI2BB2XL U1352 ( .B0(n1950), .B1(n2168), .A0N(\register[5][20] ), .A1N(
        n2169), .Y(n934) );
  OAI2BB2XL U1353 ( .B0(n1947), .B1(n2168), .A0N(\register[5][21] ), .A1N(
        n2168), .Y(n935) );
  OAI2BB2XL U1354 ( .B0(n1941), .B1(n2168), .A0N(\register[5][23] ), .A1N(
        n2168), .Y(n937) );
  OAI2BB2XL U1355 ( .B0(n1953), .B1(n2164), .A0N(\register[4][19] ), .A1N(
        n2165), .Y(n965) );
  OAI2BB2XL U1356 ( .B0(n1944), .B1(n2164), .A0N(\register[4][22] ), .A1N(
        n2164), .Y(n968) );
  OAI2BB2XL U1357 ( .B0(n1941), .B1(n2164), .A0N(\register[4][23] ), .A1N(
        n2164), .Y(n969) );
  OAI2BB2XL U1358 ( .B0(n1938), .B1(n2164), .A0N(\register[4][24] ), .A1N(
        n2164), .Y(n970) );
  OAI2BB2XL U1359 ( .B0(n1959), .B1(n2160), .A0N(\register[3][17] ), .A1N(
        n2161), .Y(n995) );
  OAI2BB2XL U1360 ( .B0(n1953), .B1(n2160), .A0N(\register[3][19] ), .A1N(
        n2161), .Y(n997) );
  OAI2BB2XL U1361 ( .B0(n1950), .B1(n2160), .A0N(\register[3][20] ), .A1N(
        n2161), .Y(n998) );
  OAI2BB2XL U1362 ( .B0(n1947), .B1(n2160), .A0N(\register[3][21] ), .A1N(
        n2160), .Y(n999) );
  OAI2BB2XL U1363 ( .B0(n1944), .B1(n2160), .A0N(\register[3][22] ), .A1N(
        n2160), .Y(n1000) );
  OAI2BB2XL U1364 ( .B0(n1941), .B1(n2160), .A0N(\register[3][23] ), .A1N(
        n2160), .Y(n1001) );
  OAI2BB2XL U1365 ( .B0(n1938), .B1(n2160), .A0N(\register[3][24] ), .A1N(
        n2160), .Y(n1002) );
  OAI2BB2XL U1366 ( .B0(n1945), .B1(n2236), .A0N(\register[22][22] ), .A1N(
        n2236), .Y(n392) );
  OAI2BB2XL U1367 ( .B0(n1942), .B1(n2236), .A0N(\register[22][23] ), .A1N(
        n2236), .Y(n393) );
  OAI2BB2XL U1368 ( .B0(n1939), .B1(n2236), .A0N(\register[22][24] ), .A1N(
        n2236), .Y(n394) );
  OAI2BB2XL U1369 ( .B0(n1960), .B1(n2228), .A0N(\register[20][17] ), .A1N(
        n2229), .Y(n451) );
  OAI2BB2XL U1370 ( .B0(n1939), .B1(n2228), .A0N(\register[20][24] ), .A1N(
        n2228), .Y(n458) );
  OAI2BB2XL U1371 ( .B0(n1954), .B1(n2220), .A0N(\register[18][19] ), .A1N(
        n2221), .Y(n517) );
  OAI2BB2XL U1372 ( .B0(n1951), .B1(n2220), .A0N(\register[18][20] ), .A1N(
        n2221), .Y(n518) );
  OAI2BB2XL U1373 ( .B0(n1948), .B1(n2220), .A0N(\register[18][21] ), .A1N(
        n2220), .Y(n519) );
  OAI2BB2XL U1374 ( .B0(n1945), .B1(n2220), .A0N(\register[18][22] ), .A1N(
        n2220), .Y(n520) );
  OAI2BB2XL U1375 ( .B0(n1942), .B1(n2220), .A0N(\register[18][23] ), .A1N(
        n2220), .Y(n521) );
  OAI2BB2XL U1376 ( .B0(n1939), .B1(n2220), .A0N(\register[18][24] ), .A1N(
        n2220), .Y(n522) );
  OAI2BB2XL U1377 ( .B0(n1963), .B1(n2212), .A0N(\register[16][16] ), .A1N(
        n2213), .Y(n578) );
  OAI2BB2XL U1378 ( .B0(n1954), .B1(n2212), .A0N(\register[16][19] ), .A1N(
        n2213), .Y(n581) );
  OAI2BB2XL U1379 ( .B0(n1951), .B1(n2212), .A0N(\register[16][20] ), .A1N(
        n2213), .Y(n582) );
  OAI2BB2XL U1380 ( .B0(n1948), .B1(n2212), .A0N(\register[16][21] ), .A1N(
        n2212), .Y(n583) );
  OAI2BB2XL U1381 ( .B0(n1945), .B1(n2212), .A0N(\register[16][22] ), .A1N(
        n2212), .Y(n584) );
  OAI2BB2XL U1382 ( .B0(n1942), .B1(n2212), .A0N(\register[16][23] ), .A1N(
        n2212), .Y(n585) );
  OAI2BB2XL U1383 ( .B0(n1939), .B1(n2212), .A0N(\register[16][24] ), .A1N(
        n2212), .Y(n586) );
  OAI2BB2XL U1384 ( .B0(n2002), .B1(n2206), .A0N(\register[15][3] ), .A1N(
        n2209), .Y(n597) );
  OAI2BB2XL U1385 ( .B0(n1999), .B1(n2206), .A0N(\register[15][4] ), .A1N(
        n2209), .Y(n598) );
  OAI2BB2XL U1386 ( .B0(n1996), .B1(n2206), .A0N(\register[15][5] ), .A1N(
        n2209), .Y(n599) );
  OAI2BB2XL U1387 ( .B0(n1993), .B1(n2206), .A0N(\register[15][6] ), .A1N(
        n2209), .Y(n600) );
  OAI2BB2XL U1388 ( .B0(n1990), .B1(n2206), .A0N(\register[15][7] ), .A1N(
        n2209), .Y(n601) );
  OAI2BB2XL U1389 ( .B0(n1987), .B1(n2207), .A0N(\register[15][8] ), .A1N(
        n2209), .Y(n602) );
  OAI2BB2XL U1390 ( .B0(n1984), .B1(n2207), .A0N(\register[15][9] ), .A1N(
        n2209), .Y(n603) );
  OAI2BB2XL U1391 ( .B0(n1981), .B1(n2207), .A0N(\register[15][10] ), .A1N(
        n2209), .Y(n604) );
  OAI2BB2XL U1392 ( .B0(n1978), .B1(n2207), .A0N(\register[15][11] ), .A1N(
        n2209), .Y(n605) );
  OAI2BB2XL U1393 ( .B0(n1975), .B1(n2207), .A0N(\register[15][12] ), .A1N(
        n2209), .Y(n606) );
  OAI2BB2XL U1394 ( .B0(n1972), .B1(n2207), .A0N(\register[15][13] ), .A1N(
        n2209), .Y(n607) );
  OAI2BB2XL U1395 ( .B0(n1969), .B1(n2207), .A0N(\register[15][14] ), .A1N(
        n2209), .Y(n608) );
  OAI2BB2XL U1396 ( .B0(n1966), .B1(n2207), .A0N(\register[15][15] ), .A1N(
        n2209), .Y(n609) );
  OAI2BB2XL U1397 ( .B0(n2005), .B1(n2202), .A0N(\register[14][2] ), .A1N(
        n2205), .Y(n628) );
  OAI2BB2XL U1398 ( .B0(n1984), .B1(n2199), .A0N(\register[13][9] ), .A1N(
        n2201), .Y(n667) );
  OAI2BB2XL U1399 ( .B0(n1992), .B1(n2190), .A0N(\register[11][6] ), .A1N(
        n2193), .Y(n728) );
  OAI2BB2XL U1400 ( .B0(n1995), .B1(n2186), .A0N(\register[10][5] ), .A1N(
        n2189), .Y(n759) );
  OAI2BB2XL U1401 ( .B0(n1992), .B1(n2186), .A0N(\register[10][6] ), .A1N(
        n2189), .Y(n760) );
  OAI2BB2XL U1402 ( .B0(n1989), .B1(n2186), .A0N(\register[10][7] ), .A1N(
        n2189), .Y(n761) );
  OAI2BB2XL U1403 ( .B0(n1986), .B1(n2187), .A0N(\register[10][8] ), .A1N(
        n2189), .Y(n762) );
  OAI2BB2XL U1404 ( .B0(n1983), .B1(n2187), .A0N(\register[10][9] ), .A1N(
        n2189), .Y(n763) );
  OAI2BB2XL U1405 ( .B0(n1980), .B1(n2187), .A0N(\register[10][10] ), .A1N(
        n2189), .Y(n764) );
  OAI2BB2XL U1406 ( .B0(n1977), .B1(n2187), .A0N(\register[10][11] ), .A1N(
        n2189), .Y(n765) );
  OAI2BB2XL U1407 ( .B0(n1974), .B1(n2187), .A0N(\register[10][12] ), .A1N(
        n2189), .Y(n766) );
  OAI2BB2XL U1408 ( .B0(n1971), .B1(n2187), .A0N(\register[10][13] ), .A1N(
        n2189), .Y(n767) );
  OAI2BB2XL U1409 ( .B0(n1968), .B1(n2187), .A0N(\register[10][14] ), .A1N(
        n2189), .Y(n768) );
  OAI2BB2XL U1410 ( .B0(n1965), .B1(n2187), .A0N(\register[10][15] ), .A1N(
        n2189), .Y(n769) );
  OAI2BB2XL U1411 ( .B0(n1962), .B1(n2188), .A0N(\register[10][16] ), .A1N(
        n2189), .Y(n770) );
  OAI2BB2XL U1412 ( .B0(n1959), .B1(n2188), .A0N(\register[10][17] ), .A1N(
        n2189), .Y(n771) );
  OAI2BB2XL U1413 ( .B0(n1956), .B1(n2187), .A0N(\register[10][18] ), .A1N(
        n2189), .Y(n772) );
  OAI2BB2XL U1414 ( .B0(n1953), .B1(n2188), .A0N(\register[10][19] ), .A1N(
        n2189), .Y(n773) );
  OAI2BB2XL U1415 ( .B0(n1935), .B1(n2187), .A0N(\register[10][25] ), .A1N(
        n2188), .Y(n779) );
  OAI2BB2XL U1416 ( .B0(n1932), .B1(n2187), .A0N(\register[10][26] ), .A1N(
        n2188), .Y(n780) );
  OAI2BB2XL U1417 ( .B0(n1929), .B1(n2187), .A0N(\register[10][27] ), .A1N(
        n2188), .Y(n781) );
  OAI2BB2XL U1418 ( .B0(n1926), .B1(n2186), .A0N(\register[10][28] ), .A1N(
        n2188), .Y(n782) );
  OAI2BB2XL U1419 ( .B0(n1920), .B1(n2186), .A0N(\register[10][30] ), .A1N(
        n2188), .Y(n784) );
  OAI2BB2XL U1420 ( .B0(n1917), .B1(n2186), .A0N(\register[10][31] ), .A1N(
        n2188), .Y(n785) );
  OAI2BB2XL U1421 ( .B0(n1935), .B1(n2183), .A0N(\register[9][25] ), .A1N(
        n2184), .Y(n811) );
  OAI2BB2XL U1422 ( .B0(n1932), .B1(n2183), .A0N(\register[9][26] ), .A1N(
        n2184), .Y(n812) );
  OAI2BB2XL U1423 ( .B0(n1926), .B1(n2182), .A0N(\register[9][28] ), .A1N(
        n2184), .Y(n814) );
  OAI2BB2XL U1424 ( .B0(n1923), .B1(n2182), .A0N(\register[9][29] ), .A1N(
        n2184), .Y(n815) );
  OAI2BB2XL U1425 ( .B0(n1920), .B1(n2182), .A0N(\register[9][30] ), .A1N(
        n2184), .Y(n816) );
  OAI2BB2XL U1426 ( .B0(n1935), .B1(n2179), .A0N(\register[8][25] ), .A1N(
        n2180), .Y(n843) );
  OAI2BB2XL U1427 ( .B0(n1932), .B1(n2179), .A0N(\register[8][26] ), .A1N(
        n2180), .Y(n844) );
  OAI2BB2XL U1428 ( .B0(n1929), .B1(n2179), .A0N(\register[8][27] ), .A1N(
        n2180), .Y(n845) );
  OAI2BB2XL U1429 ( .B0(n1926), .B1(n2178), .A0N(\register[8][28] ), .A1N(
        n2180), .Y(n846) );
  OAI2BB2XL U1430 ( .B0(n1920), .B1(n2178), .A0N(\register[8][30] ), .A1N(
        n2180), .Y(n848) );
  OAI2BB2XL U1431 ( .B0(n1968), .B1(n2175), .A0N(\register[7][14] ), .A1N(
        n2177), .Y(n864) );
  OAI2BB2XL U1432 ( .B0(n1959), .B1(n2176), .A0N(\register[7][17] ), .A1N(
        n2177), .Y(n867) );
  OAI2BB2XL U1433 ( .B0(n1944), .B1(n2176), .A0N(\register[7][22] ), .A1N(
        n2176), .Y(n872) );
  OAI2BB2XL U1434 ( .B0(n1941), .B1(n2176), .A0N(\register[7][23] ), .A1N(
        n2176), .Y(n873) );
  OAI2BB2XL U1435 ( .B0(n1938), .B1(n2176), .A0N(\register[7][24] ), .A1N(
        n2176), .Y(n874) );
  OAI2BB2XL U1436 ( .B0(n1941), .B1(n2172), .A0N(\register[6][23] ), .A1N(
        n2172), .Y(n905) );
  OAI2BB2XL U1437 ( .B0(n1944), .B1(n2168), .A0N(\register[5][22] ), .A1N(
        n2168), .Y(n936) );
  OAI2BB2XL U1438 ( .B0(n1935), .B1(n2167), .A0N(\register[5][25] ), .A1N(
        n2168), .Y(n939) );
  OAI2BB2XL U1439 ( .B0(n1932), .B1(n2167), .A0N(\register[5][26] ), .A1N(
        n2168), .Y(n940) );
  OAI2BB2XL U1440 ( .B0(n1929), .B1(n2167), .A0N(\register[5][27] ), .A1N(
        n2168), .Y(n941) );
  OAI2BB2XL U1441 ( .B0(n1926), .B1(n2166), .A0N(\register[5][28] ), .A1N(
        n2168), .Y(n942) );
  OAI2BB2XL U1442 ( .B0(n1920), .B1(n2166), .A0N(\register[5][30] ), .A1N(
        n2168), .Y(n944) );
  OAI2BB2XL U1443 ( .B0(n2010), .B1(n2162), .A0N(\register[4][0] ), .A1N(n2164), .Y(n946) );
  OAI2BB2XL U1444 ( .B0(n2007), .B1(n2162), .A0N(\register[4][1] ), .A1N(n2165), .Y(n947) );
  OAI2BB2XL U1445 ( .B0(n2004), .B1(n2162), .A0N(\register[4][2] ), .A1N(n2165), .Y(n948) );
  OAI2BB2XL U1446 ( .B0(n2001), .B1(n2162), .A0N(\register[4][3] ), .A1N(n2165), .Y(n949) );
  OAI2BB2XL U1447 ( .B0(n1989), .B1(n2162), .A0N(\register[4][7] ), .A1N(n2165), .Y(n953) );
  OAI2BB2XL U1448 ( .B0(n1986), .B1(n2163), .A0N(\register[4][8] ), .A1N(n2165), .Y(n954) );
  OAI2BB2XL U1449 ( .B0(n1983), .B1(n2163), .A0N(\register[4][9] ), .A1N(n2165), .Y(n955) );
  OAI2BB2XL U1450 ( .B0(n1980), .B1(n2163), .A0N(\register[4][10] ), .A1N(
        n2165), .Y(n956) );
  OAI2BB2XL U1451 ( .B0(n1977), .B1(n2163), .A0N(\register[4][11] ), .A1N(
        n2165), .Y(n957) );
  OAI2BB2XL U1452 ( .B0(n1974), .B1(n2163), .A0N(\register[4][12] ), .A1N(
        n2165), .Y(n958) );
  OAI2BB2XL U1453 ( .B0(n1965), .B1(n2163), .A0N(\register[4][15] ), .A1N(
        n2165), .Y(n961) );
  OAI2BB2XL U1454 ( .B0(n1962), .B1(n2164), .A0N(\register[4][16] ), .A1N(
        n2165), .Y(n962) );
  OAI2BB2XL U1455 ( .B0(n1959), .B1(n2164), .A0N(\register[4][17] ), .A1N(
        n2165), .Y(n963) );
  OAI2BB2XL U1456 ( .B0(n1956), .B1(n2163), .A0N(\register[4][18] ), .A1N(
        n2165), .Y(n964) );
  OAI2BB2XL U1457 ( .B0(n1950), .B1(n2164), .A0N(\register[4][20] ), .A1N(
        n2165), .Y(n966) );
  OAI2BB2XL U1458 ( .B0(n1947), .B1(n2164), .A0N(\register[4][21] ), .A1N(
        n2164), .Y(n967) );
  OAI2BB2XL U1459 ( .B0(n1960), .B1(n2212), .A0N(\register[16][17] ), .A1N(
        n2213), .Y(n579) );
  OAI2BB2XL U1460 ( .B0(n1956), .B1(n2175), .A0N(\register[7][18] ), .A1N(
        n2177), .Y(n868) );
  OAI2BB2XL U1461 ( .B0(n1935), .B1(n2175), .A0N(\register[7][25] ), .A1N(
        n2176), .Y(n875) );
  OAI2BB2XL U1462 ( .B0(n1932), .B1(n2175), .A0N(\register[7][26] ), .A1N(
        n2176), .Y(n876) );
  OAI2BB2XL U1463 ( .B0(n1935), .B1(n2163), .A0N(\register[4][25] ), .A1N(
        n2164), .Y(n971) );
  OAI2BB2XL U1464 ( .B0(n1929), .B1(n2163), .A0N(\register[4][27] ), .A1N(
        n2164), .Y(n973) );
  OAI2BB2XL U1465 ( .B0(n1926), .B1(n2162), .A0N(\register[4][28] ), .A1N(
        n2164), .Y(n974) );
  OAI2BB2XL U1466 ( .B0(n1920), .B1(n2162), .A0N(\register[4][30] ), .A1N(
        n2164), .Y(n976) );
  OAI2BB2XL U1467 ( .B0(n1917), .B1(n2162), .A0N(\register[4][31] ), .A1N(
        n2164), .Y(n977) );
  OAI2BB2XL U1468 ( .B0(n2010), .B1(n2158), .A0N(\register[3][0] ), .A1N(n2160), .Y(n978) );
  OAI2BB2XL U1469 ( .B0(n2007), .B1(n2158), .A0N(\register[3][1] ), .A1N(n2161), .Y(n979) );
  OAI2BB2XL U1470 ( .B0(n1998), .B1(n2158), .A0N(\register[3][4] ), .A1N(n2161), .Y(n982) );
  OAI2BB2XL U1471 ( .B0(n1995), .B1(n2158), .A0N(\register[3][5] ), .A1N(n2161), .Y(n983) );
  OAI2BB2XL U1472 ( .B0(n1992), .B1(n2158), .A0N(\register[3][6] ), .A1N(n2161), .Y(n984) );
  OAI2BB2XL U1473 ( .B0(n1989), .B1(n2158), .A0N(\register[3][7] ), .A1N(n2161), .Y(n985) );
  OAI2BB2XL U1474 ( .B0(n1986), .B1(n2159), .A0N(\register[3][8] ), .A1N(n2161), .Y(n986) );
  OAI2BB2XL U1475 ( .B0(n1983), .B1(n2159), .A0N(\register[3][9] ), .A1N(n2161), .Y(n987) );
  OAI2BB2XL U1476 ( .B0(n1980), .B1(n2159), .A0N(\register[3][10] ), .A1N(
        n2161), .Y(n988) );
  OAI2BB2XL U1477 ( .B0(n1977), .B1(n2159), .A0N(\register[3][11] ), .A1N(
        n2161), .Y(n989) );
  OAI2BB2XL U1478 ( .B0(n1971), .B1(n2159), .A0N(\register[3][13] ), .A1N(
        n2161), .Y(n991) );
  OAI2BB2XL U1479 ( .B0(n1968), .B1(n2159), .A0N(\register[3][14] ), .A1N(
        n2161), .Y(n992) );
  OAI2BB2XL U1480 ( .B0(n1965), .B1(n2159), .A0N(\register[3][15] ), .A1N(
        n2161), .Y(n993) );
  OAI2BB2XL U1481 ( .B0(n1962), .B1(n2160), .A0N(\register[3][16] ), .A1N(
        n2161), .Y(n994) );
  OAI2BB2XL U1482 ( .B0(n1956), .B1(n2159), .A0N(\register[3][18] ), .A1N(
        n2161), .Y(n996) );
  OAI2BB2XL U1483 ( .B0(n1935), .B1(n2159), .A0N(\register[3][25] ), .A1N(
        n2160), .Y(n1003) );
  OAI2BB2XL U1484 ( .B0(n1932), .B1(n2159), .A0N(\register[3][26] ), .A1N(
        n2160), .Y(n1004) );
  OAI2BB2XL U1485 ( .B0(n1929), .B1(n2159), .A0N(\register[3][27] ), .A1N(
        n2160), .Y(n1005) );
  OAI2BB2XL U1486 ( .B0(n1926), .B1(n2158), .A0N(\register[3][28] ), .A1N(
        n2160), .Y(n1006) );
  OAI2BB2XL U1487 ( .B0(n1923), .B1(n2158), .A0N(\register[3][29] ), .A1N(
        n2160), .Y(n1007) );
  OAI2BB2XL U1488 ( .B0(n1920), .B1(n2158), .A0N(\register[3][30] ), .A1N(
        n2160), .Y(n1008) );
  OAI2BB2XL U1489 ( .B0(n1917), .B1(n2158), .A0N(\register[3][31] ), .A1N(
        n2160), .Y(n1009) );
  OAI2BB2XL U1490 ( .B0(n2010), .B1(n2154), .A0N(\register[2][0] ), .A1N(n2156), .Y(n1010) );
  OAI2BB2XL U1491 ( .B0(n2007), .B1(n2154), .A0N(\register[2][1] ), .A1N(n2157), .Y(n1011) );
  OAI2BB2XL U1492 ( .B0(n2004), .B1(n2154), .A0N(\register[2][2] ), .A1N(n2157), .Y(n1012) );
  OAI2BB2XL U1493 ( .B0(n2001), .B1(n2154), .A0N(\register[2][3] ), .A1N(n2157), .Y(n1013) );
  OAI2BB2XL U1494 ( .B0(n1998), .B1(n2154), .A0N(\register[2][4] ), .A1N(n2157), .Y(n1014) );
  OAI2BB2XL U1495 ( .B0(n1995), .B1(n2154), .A0N(\register[2][5] ), .A1N(n2157), .Y(n1015) );
  OAI2BB2XL U1496 ( .B0(n1992), .B1(n2154), .A0N(\register[2][6] ), .A1N(n2157), .Y(n1016) );
  OAI2BB2XL U1497 ( .B0(n1989), .B1(n2154), .A0N(\register[2][7] ), .A1N(n2157), .Y(n1017) );
  OAI2BB2XL U1498 ( .B0(n1986), .B1(n2155), .A0N(\register[2][8] ), .A1N(n2157), .Y(n1018) );
  OAI2BB2XL U1499 ( .B0(n1983), .B1(n2155), .A0N(\register[2][9] ), .A1N(n2157), .Y(n1019) );
  OAI2BB2XL U1500 ( .B0(n1980), .B1(n2155), .A0N(\register[2][10] ), .A1N(
        n2157), .Y(n1020) );
  OAI2BB2XL U1501 ( .B0(n1977), .B1(n2155), .A0N(\register[2][11] ), .A1N(
        n2157), .Y(n1021) );
  OAI2BB2XL U1502 ( .B0(n1974), .B1(n2155), .A0N(\register[2][12] ), .A1N(
        n2157), .Y(n1022) );
  OAI2BB2XL U1503 ( .B0(n1971), .B1(n2155), .A0N(\register[2][13] ), .A1N(
        n2157), .Y(n1023) );
  OAI2BB2XL U1504 ( .B0(n1965), .B1(n2155), .A0N(\register[2][15] ), .A1N(
        n2157), .Y(n1025) );
  OAI2BB2XL U1505 ( .B0(n1962), .B1(n2156), .A0N(\register[2][16] ), .A1N(
        n2157), .Y(n1026) );
  OAI2BB2XL U1506 ( .B0(n1959), .B1(n2156), .A0N(\register[2][17] ), .A1N(
        n2157), .Y(n1027) );
  OAI2BB2XL U1507 ( .B0(n1956), .B1(n2155), .A0N(\register[2][18] ), .A1N(
        n2157), .Y(n1028) );
  OAI2BB2XL U1508 ( .B0(n1953), .B1(n2156), .A0N(\register[2][19] ), .A1N(
        n2157), .Y(n1029) );
  OAI2BB2XL U1509 ( .B0(n1950), .B1(n2156), .A0N(\register[2][20] ), .A1N(
        n2157), .Y(n1030) );
  OAI2BB2XL U1510 ( .B0(n1947), .B1(n2156), .A0N(\register[2][21] ), .A1N(
        n2156), .Y(n1031) );
  OAI2BB2XL U1511 ( .B0(n1944), .B1(n2156), .A0N(\register[2][22] ), .A1N(
        n2156), .Y(n1032) );
  OAI2BB2XL U1512 ( .B0(n1941), .B1(n2156), .A0N(\register[2][23] ), .A1N(
        n2156), .Y(n1033) );
  OAI2BB2XL U1513 ( .B0(n1938), .B1(n2156), .A0N(\register[2][24] ), .A1N(
        n2156), .Y(n1034) );
  OAI2BB2XL U1514 ( .B0(n1935), .B1(n2155), .A0N(\register[2][25] ), .A1N(
        n2156), .Y(n1035) );
  OAI2BB2XL U1515 ( .B0(n1932), .B1(n2155), .A0N(\register[2][26] ), .A1N(
        n2156), .Y(n1036) );
  OAI2BB2XL U1516 ( .B0(n1929), .B1(n2155), .A0N(\register[2][27] ), .A1N(
        n2156), .Y(n1037) );
  OAI2BB2XL U1517 ( .B0(n1926), .B1(n2154), .A0N(\register[2][28] ), .A1N(
        n2156), .Y(n1038) );
  OAI2BB2XL U1518 ( .B0(n1923), .B1(n2154), .A0N(\register[2][29] ), .A1N(
        n2156), .Y(n1039) );
  OAI2BB2XL U1519 ( .B0(n2007), .B1(n2150), .A0N(\register[1][1] ), .A1N(n2153), .Y(n1043) );
  OAI2BB2XL U1520 ( .B0(n2004), .B1(n2150), .A0N(\register[1][2] ), .A1N(n2153), .Y(n1044) );
  OAI2BB2XL U1521 ( .B0(n1995), .B1(n2150), .A0N(\register[1][5] ), .A1N(n2153), .Y(n1047) );
  OAI2BB2XL U1522 ( .B0(n1989), .B1(n2150), .A0N(\register[1][7] ), .A1N(n2153), .Y(n1049) );
  OAI2BB2XL U1523 ( .B0(n1986), .B1(n2151), .A0N(\register[1][8] ), .A1N(n2153), .Y(n1050) );
  OAI2BB2XL U1524 ( .B0(n1983), .B1(n2151), .A0N(\register[1][9] ), .A1N(n2153), .Y(n1051) );
  OAI2BB2XL U1525 ( .B0(n1980), .B1(n2151), .A0N(\register[1][10] ), .A1N(
        n2153), .Y(n1052) );
  OAI2BB2XL U1526 ( .B0(n1974), .B1(n2151), .A0N(\register[1][12] ), .A1N(
        n2153), .Y(n1054) );
  OAI2BB2XL U1527 ( .B0(n1968), .B1(n2151), .A0N(\register[1][14] ), .A1N(
        n2153), .Y(n1056) );
  OAI2BB2XL U1528 ( .B0(n1959), .B1(n2152), .A0N(\register[1][17] ), .A1N(
        n2153), .Y(n1059) );
  OAI2BB2XL U1529 ( .B0(n1956), .B1(n2151), .A0N(\register[1][18] ), .A1N(
        n2153), .Y(n1060) );
  OAI2BB2XL U1530 ( .B0(n1953), .B1(n2152), .A0N(\register[1][19] ), .A1N(
        n2153), .Y(n1061) );
  OAI2BB2XL U1531 ( .B0(n1950), .B1(n2152), .A0N(\register[1][20] ), .A1N(
        n2153), .Y(n1062) );
  OAI2BB2XL U1532 ( .B0(n1947), .B1(n2152), .A0N(\register[1][21] ), .A1N(
        n2152), .Y(n1063) );
  OAI2BB2XL U1533 ( .B0(n1944), .B1(n2152), .A0N(\register[1][22] ), .A1N(
        n2152), .Y(n1064) );
  OAI2BB2XL U1534 ( .B0(n1941), .B1(n2152), .A0N(\register[1][23] ), .A1N(
        n2152), .Y(n1065) );
  OAI2BB2XL U1535 ( .B0(n1938), .B1(n2152), .A0N(\register[1][24] ), .A1N(
        n2152), .Y(n1066) );
  OAI2BB2XL U1536 ( .B0(n1929), .B1(n2151), .A0N(\register[1][27] ), .A1N(
        n2152), .Y(n1069) );
  OAI2BB2XL U1537 ( .B0(n1926), .B1(n2150), .A0N(\register[1][28] ), .A1N(
        n2152), .Y(n1070) );
  OAI2BB2XL U1538 ( .B0(n1923), .B1(n2150), .A0N(\register[1][29] ), .A1N(
        n2152), .Y(n1071) );
  OAI2BB2XL U1539 ( .B0(n1920), .B1(n2150), .A0N(\register[1][30] ), .A1N(
        n2152), .Y(n1072) );
  OAI2BB2XL U1540 ( .B0(n1917), .B1(n2150), .A0N(\register[1][31] ), .A1N(
        n2152), .Y(n1073) );
  OAI2BB2XL U1541 ( .B0(n2010), .B1(n2146), .A0N(\register[0][0] ), .A1N(n2148), .Y(n1074) );
  OAI2BB2XL U1542 ( .B0(n2007), .B1(n2146), .A0N(\register[0][1] ), .A1N(n2149), .Y(n1075) );
  OAI2BB2XL U1543 ( .B0(n2004), .B1(n2146), .A0N(\register[0][2] ), .A1N(n2149), .Y(n1076) );
  OAI2BB2XL U1544 ( .B0(n2001), .B1(n2146), .A0N(\register[0][3] ), .A1N(n2149), .Y(n1077) );
  OAI2BB2XL U1545 ( .B0(n1998), .B1(n2146), .A0N(\register[0][4] ), .A1N(n2149), .Y(n1078) );
  OAI2BB2XL U1546 ( .B0(n1995), .B1(n2146), .A0N(\register[0][5] ), .A1N(n2149), .Y(n1079) );
  OAI2BB2XL U1547 ( .B0(n1992), .B1(n2146), .A0N(\register[0][6] ), .A1N(n2149), .Y(n1080) );
  OAI2BB2XL U1548 ( .B0(n1989), .B1(n2146), .A0N(\register[0][7] ), .A1N(n2149), .Y(n1081) );
  OAI2BB2XL U1549 ( .B0(n1986), .B1(n2147), .A0N(\register[0][8] ), .A1N(n2149), .Y(n1082) );
  OAI2BB2XL U1550 ( .B0(n1983), .B1(n2147), .A0N(\register[0][9] ), .A1N(n2149), .Y(n1083) );
  OAI2BB2XL U1551 ( .B0(n1980), .B1(n2147), .A0N(\register[0][10] ), .A1N(
        n2149), .Y(n1084) );
  OAI2BB2XL U1552 ( .B0(n1977), .B1(n2147), .A0N(\register[0][11] ), .A1N(
        n2149), .Y(n1085) );
  OAI2BB2XL U1553 ( .B0(n1974), .B1(n2147), .A0N(\register[0][12] ), .A1N(
        n2149), .Y(n1086) );
  OAI2BB2XL U1554 ( .B0(n1971), .B1(n2147), .A0N(\register[0][13] ), .A1N(
        n2149), .Y(n1087) );
  OAI2BB2XL U1555 ( .B0(n1968), .B1(n2147), .A0N(\register[0][14] ), .A1N(
        n2149), .Y(n1088) );
  OAI2BB2XL U1556 ( .B0(n1965), .B1(n2147), .A0N(\register[0][15] ), .A1N(
        n2149), .Y(n1089) );
  OAI2BB2XL U1557 ( .B0(n1962), .B1(n2148), .A0N(\register[0][16] ), .A1N(
        n2149), .Y(n1090) );
  OAI2BB2XL U1558 ( .B0(n1959), .B1(n2148), .A0N(\register[0][17] ), .A1N(
        n2149), .Y(n1091) );
  OAI2BB2XL U1559 ( .B0(n1956), .B1(n2147), .A0N(\register[0][18] ), .A1N(
        n2149), .Y(n1092) );
  OAI2BB2XL U1560 ( .B0(n1953), .B1(n2148), .A0N(\register[0][19] ), .A1N(
        n2149), .Y(n1093) );
  OAI2BB2XL U1561 ( .B0(n1950), .B1(n2148), .A0N(\register[0][20] ), .A1N(
        n2149), .Y(n1094) );
  OAI2BB2XL U1562 ( .B0(n1947), .B1(n2148), .A0N(\register[0][21] ), .A1N(
        n2148), .Y(n1095) );
  OAI2BB2XL U1563 ( .B0(n1941), .B1(n2148), .A0N(\register[0][23] ), .A1N(
        n2148), .Y(n1097) );
  OAI2BB2XL U1564 ( .B0(n1938), .B1(n2148), .A0N(\register[0][24] ), .A1N(
        n2148), .Y(n1098) );
  OAI2BB2XL U1565 ( .B0(n2011), .B1(n2238), .A0N(\register[23][0] ), .A1N(
        n2240), .Y(n338) );
  OAI2BB2XL U1566 ( .B0(n2008), .B1(n2238), .A0N(\register[23][1] ), .A1N(
        n2241), .Y(n339) );
  OAI2BB2XL U1567 ( .B0(n2005), .B1(n2238), .A0N(\register[23][2] ), .A1N(
        n2241), .Y(n340) );
  OAI2BB2XL U1568 ( .B0(n2002), .B1(n2238), .A0N(\register[23][3] ), .A1N(
        n2241), .Y(n341) );
  OAI2BB2XL U1569 ( .B0(n1999), .B1(n2238), .A0N(\register[23][4] ), .A1N(
        n2241), .Y(n342) );
  OAI2BB2XL U1570 ( .B0(n1996), .B1(n2238), .A0N(\register[23][5] ), .A1N(
        n2241), .Y(n343) );
  OAI2BB2XL U1571 ( .B0(n1993), .B1(n2238), .A0N(\register[23][6] ), .A1N(
        n2241), .Y(n344) );
  OAI2BB2XL U1572 ( .B0(n1990), .B1(n2238), .A0N(\register[23][7] ), .A1N(
        n2241), .Y(n345) );
  OAI2BB2XL U1573 ( .B0(n1987), .B1(n2239), .A0N(\register[23][8] ), .A1N(
        n2241), .Y(n346) );
  OAI2BB2XL U1574 ( .B0(n1984), .B1(n2239), .A0N(\register[23][9] ), .A1N(
        n2241), .Y(n347) );
  OAI2BB2XL U1575 ( .B0(n1981), .B1(n2239), .A0N(\register[23][10] ), .A1N(
        n2241), .Y(n348) );
  OAI2BB2XL U1576 ( .B0(n1978), .B1(n2239), .A0N(\register[23][11] ), .A1N(
        n2241), .Y(n349) );
  OAI2BB2XL U1577 ( .B0(n1975), .B1(n2239), .A0N(\register[23][12] ), .A1N(
        n2241), .Y(n350) );
  OAI2BB2XL U1578 ( .B0(n1972), .B1(n2239), .A0N(\register[23][13] ), .A1N(
        n2241), .Y(n351) );
  OAI2BB2XL U1579 ( .B0(n1969), .B1(n2239), .A0N(\register[23][14] ), .A1N(
        n2241), .Y(n352) );
  OAI2BB2XL U1580 ( .B0(n1966), .B1(n2239), .A0N(\register[23][15] ), .A1N(
        n2241), .Y(n353) );
  OAI2BB2XL U1581 ( .B0(n1963), .B1(n2240), .A0N(\register[23][16] ), .A1N(
        n2241), .Y(n354) );
  OAI2BB2XL U1582 ( .B0(n1960), .B1(n2240), .A0N(\register[23][17] ), .A1N(
        n2241), .Y(n355) );
  OAI2BB2XL U1583 ( .B0(n1954), .B1(n2240), .A0N(\register[23][19] ), .A1N(
        n2241), .Y(n357) );
  OAI2BB2XL U1584 ( .B0(n1951), .B1(n2240), .A0N(\register[23][20] ), .A1N(
        n2241), .Y(n358) );
  OAI2BB2XL U1585 ( .B0(n1948), .B1(n2240), .A0N(\register[23][21] ), .A1N(
        n2240), .Y(n359) );
  OAI2BB2XL U1586 ( .B0(n1939), .B1(n2240), .A0N(\register[23][24] ), .A1N(
        n2240), .Y(n362) );
  OAI2BB2XL U1587 ( .B0(n1918), .B1(n2238), .A0N(\register[23][31] ), .A1N(
        n2240), .Y(n369) );
  OAI2BB2XL U1588 ( .B0(n2011), .B1(n2234), .A0N(\register[22][0] ), .A1N(
        n2236), .Y(n370) );
  OAI2BB2XL U1589 ( .B0(n2008), .B1(n2234), .A0N(\register[22][1] ), .A1N(
        n2237), .Y(n371) );
  OAI2BB2XL U1590 ( .B0(n2005), .B1(n2234), .A0N(\register[22][2] ), .A1N(
        n2237), .Y(n372) );
  OAI2BB2XL U1591 ( .B0(n2002), .B1(n2234), .A0N(\register[22][3] ), .A1N(
        n2237), .Y(n373) );
  OAI2BB2XL U1592 ( .B0(n1999), .B1(n2234), .A0N(\register[22][4] ), .A1N(
        n2237), .Y(n374) );
  OAI2BB2XL U1593 ( .B0(n1996), .B1(n2234), .A0N(\register[22][5] ), .A1N(
        n2237), .Y(n375) );
  OAI2BB2XL U1594 ( .B0(n1993), .B1(n2234), .A0N(\register[22][6] ), .A1N(
        n2237), .Y(n376) );
  OAI2BB2XL U1595 ( .B0(n1990), .B1(n2234), .A0N(\register[22][7] ), .A1N(
        n2237), .Y(n377) );
  OAI2BB2XL U1596 ( .B0(n1987), .B1(n2235), .A0N(\register[22][8] ), .A1N(
        n2237), .Y(n378) );
  OAI2BB2XL U1597 ( .B0(n1984), .B1(n2235), .A0N(\register[22][9] ), .A1N(
        n2237), .Y(n379) );
  OAI2BB2XL U1598 ( .B0(n1981), .B1(n2235), .A0N(\register[22][10] ), .A1N(
        n2237), .Y(n380) );
  OAI2BB2XL U1599 ( .B0(n1978), .B1(n2235), .A0N(\register[22][11] ), .A1N(
        n2237), .Y(n381) );
  OAI2BB2XL U1600 ( .B0(n1975), .B1(n2235), .A0N(\register[22][12] ), .A1N(
        n2237), .Y(n382) );
  OAI2BB2XL U1601 ( .B0(n1972), .B1(n2235), .A0N(\register[22][13] ), .A1N(
        n2237), .Y(n383) );
  OAI2BB2XL U1602 ( .B0(n1969), .B1(n2235), .A0N(\register[22][14] ), .A1N(
        n2237), .Y(n384) );
  OAI2BB2XL U1603 ( .B0(n1966), .B1(n2235), .A0N(\register[22][15] ), .A1N(
        n2237), .Y(n385) );
  OAI2BB2XL U1604 ( .B0(n1963), .B1(n2236), .A0N(\register[22][16] ), .A1N(
        n2237), .Y(n386) );
  OAI2BB2XL U1605 ( .B0(n1960), .B1(n2236), .A0N(\register[22][17] ), .A1N(
        n2237), .Y(n387) );
  OAI2BB2XL U1606 ( .B0(n1954), .B1(n2236), .A0N(\register[22][19] ), .A1N(
        n2237), .Y(n389) );
  OAI2BB2XL U1607 ( .B0(n1951), .B1(n2236), .A0N(\register[22][20] ), .A1N(
        n2237), .Y(n390) );
  OAI2BB2XL U1608 ( .B0(n1948), .B1(n2236), .A0N(\register[22][21] ), .A1N(
        n2236), .Y(n391) );
  OAI2BB2XL U1609 ( .B0(n1954), .B1(n2224), .A0N(\register[19][19] ), .A1N(
        n2225), .Y(n485) );
  OAI2BB2XL U1610 ( .B0(n1989), .B1(n2190), .A0N(\register[11][7] ), .A1N(
        n2193), .Y(n729) );
  OAI2BB2XL U1611 ( .B0(n1986), .B1(n2191), .A0N(\register[11][8] ), .A1N(
        n2193), .Y(n730) );
  OAI2BB2XL U1612 ( .B0(n1917), .B1(n2190), .A0N(\register[11][31] ), .A1N(
        n2192), .Y(n753) );
  OAI2BB2XL U1613 ( .B0(n2010), .B1(n2186), .A0N(\register[10][0] ), .A1N(
        n2188), .Y(n754) );
  OAI2BB2XL U1614 ( .B0(n2007), .B1(n2186), .A0N(\register[10][1] ), .A1N(
        n2189), .Y(n755) );
  OAI2BB2XL U1615 ( .B0(n2004), .B1(n2186), .A0N(\register[10][2] ), .A1N(
        n2189), .Y(n756) );
  OAI2BB2XL U1616 ( .B0(n2001), .B1(n2186), .A0N(\register[10][3] ), .A1N(
        n2189), .Y(n757) );
  OAI2BB2XL U1617 ( .B0(n1998), .B1(n2186), .A0N(\register[10][4] ), .A1N(
        n2189), .Y(n758) );
  OAI2BB2XL U1618 ( .B0(n1938), .B1(n2168), .A0N(\register[5][24] ), .A1N(
        n2168), .Y(n938) );
  OAI2BB2XL U1619 ( .B0(n1923), .B1(n2166), .A0N(\register[5][29] ), .A1N(
        n2168), .Y(n943) );
  OAI2BB2XL U1620 ( .B0(n1917), .B1(n2166), .A0N(\register[5][31] ), .A1N(
        n2168), .Y(n945) );
  OAI2BB2XL U1621 ( .B0(n1998), .B1(n2162), .A0N(\register[4][4] ), .A1N(n2165), .Y(n950) );
  OAI2BB2XL U1622 ( .B0(n1995), .B1(n2162), .A0N(\register[4][5] ), .A1N(n2165), .Y(n951) );
  OAI2BB2XL U1623 ( .B0(n1971), .B1(n2163), .A0N(\register[4][13] ), .A1N(
        n2165), .Y(n959) );
  OAI2BB2XL U1624 ( .B0(n1917), .B1(n2154), .A0N(\register[2][31] ), .A1N(
        n2156), .Y(n1041) );
  OAI2BB2XL U1625 ( .B0(n2010), .B1(n2150), .A0N(\register[1][0] ), .A1N(n2152), .Y(n1042) );
  OAI2BB2XL U1626 ( .B0(n2001), .B1(n2150), .A0N(\register[1][3] ), .A1N(n2153), .Y(n1045) );
  OAI2BB2XL U1627 ( .B0(n1998), .B1(n2150), .A0N(\register[1][4] ), .A1N(n2153), .Y(n1046) );
  OAI2BB2XL U1628 ( .B0(n1944), .B1(n2148), .A0N(\register[0][22] ), .A1N(
        n2148), .Y(n1096) );
  OAI2BB2XL U1629 ( .B0(n1935), .B1(n2147), .A0N(\register[0][25] ), .A1N(
        n2148), .Y(n1099) );
  OAI2BB2XL U1630 ( .B0(n1926), .B1(n2146), .A0N(\register[0][28] ), .A1N(
        n2148), .Y(n1102) );
  OAI2BB2XL U1631 ( .B0(n1923), .B1(n2146), .A0N(\register[0][29] ), .A1N(
        n2148), .Y(n1103) );
  OAI2BB2XL U1632 ( .B0(n1957), .B1(n2239), .A0N(\register[23][18] ), .A1N(
        n2241), .Y(n356) );
  OAI2BB2XL U1633 ( .B0(n1945), .B1(n2240), .A0N(\register[23][22] ), .A1N(
        n2240), .Y(n360) );
  OAI2BB2XL U1634 ( .B0(n1942), .B1(n2240), .A0N(\register[23][23] ), .A1N(
        n2240), .Y(n361) );
  OAI2BB2XL U1635 ( .B0(n1936), .B1(n2239), .A0N(\register[23][25] ), .A1N(
        n2240), .Y(n363) );
  OAI2BB2XL U1636 ( .B0(n1933), .B1(n2239), .A0N(\register[23][26] ), .A1N(
        n2240), .Y(n364) );
  OAI2BB2XL U1637 ( .B0(n1930), .B1(n2239), .A0N(\register[23][27] ), .A1N(
        n2240), .Y(n365) );
  OAI2BB2XL U1638 ( .B0(n1927), .B1(n2238), .A0N(\register[23][28] ), .A1N(
        n2240), .Y(n366) );
  OAI2BB2XL U1639 ( .B0(n1924), .B1(n2238), .A0N(\register[23][29] ), .A1N(
        n2240), .Y(n367) );
  OAI2BB2XL U1640 ( .B0(n1921), .B1(n2238), .A0N(\register[23][30] ), .A1N(
        n2240), .Y(n368) );
  OAI2BB2XL U1641 ( .B0(n1957), .B1(n2235), .A0N(\register[22][18] ), .A1N(
        n2237), .Y(n388) );
  OAI2BB2XL U1642 ( .B0(n1936), .B1(n2235), .A0N(\register[22][25] ), .A1N(
        n2236), .Y(n395) );
  OAI2BB2XL U1643 ( .B0(n1933), .B1(n2235), .A0N(\register[22][26] ), .A1N(
        n2236), .Y(n396) );
  OAI2BB2XL U1644 ( .B0(n1930), .B1(n2235), .A0N(\register[22][27] ), .A1N(
        n2236), .Y(n397) );
  OAI2BB2XL U1645 ( .B0(n1927), .B1(n2234), .A0N(\register[22][28] ), .A1N(
        n2236), .Y(n398) );
  OAI2BB2XL U1646 ( .B0(n1924), .B1(n2234), .A0N(\register[22][29] ), .A1N(
        n2236), .Y(n399) );
  OAI2BB2XL U1647 ( .B0(n1921), .B1(n2234), .A0N(\register[22][30] ), .A1N(
        n2236), .Y(n400) );
  OAI2BB2XL U1648 ( .B0(n1918), .B1(n2234), .A0N(\register[22][31] ), .A1N(
        n2236), .Y(n401) );
  OAI2BB2XL U1649 ( .B0(n2011), .B1(n2230), .A0N(\register[21][0] ), .A1N(
        n2232), .Y(n402) );
  OAI2BB2XL U1650 ( .B0(n2008), .B1(n2230), .A0N(\register[21][1] ), .A1N(
        n2233), .Y(n403) );
  OAI2BB2XL U1651 ( .B0(n2005), .B1(n2230), .A0N(\register[21][2] ), .A1N(
        n2233), .Y(n404) );
  OAI2BB2XL U1652 ( .B0(n2002), .B1(n2230), .A0N(\register[21][3] ), .A1N(
        n2233), .Y(n405) );
  OAI2BB2XL U1653 ( .B0(n1999), .B1(n2230), .A0N(\register[21][4] ), .A1N(
        n2233), .Y(n406) );
  OAI2BB2XL U1654 ( .B0(n1996), .B1(n2230), .A0N(\register[21][5] ), .A1N(
        n2233), .Y(n407) );
  OAI2BB2XL U1655 ( .B0(n1993), .B1(n2230), .A0N(\register[21][6] ), .A1N(
        n2233), .Y(n408) );
  OAI2BB2XL U1656 ( .B0(n1990), .B1(n2230), .A0N(\register[21][7] ), .A1N(
        n2233), .Y(n409) );
  OAI2BB2XL U1657 ( .B0(n1987), .B1(n2231), .A0N(\register[21][8] ), .A1N(
        n2233), .Y(n410) );
  OAI2BB2XL U1658 ( .B0(n1984), .B1(n2231), .A0N(\register[21][9] ), .A1N(
        n2233), .Y(n411) );
  OAI2BB2XL U1659 ( .B0(n1981), .B1(n2231), .A0N(\register[21][10] ), .A1N(
        n2233), .Y(n412) );
  OAI2BB2XL U1660 ( .B0(n1978), .B1(n2231), .A0N(\register[21][11] ), .A1N(
        n2233), .Y(n413) );
  OAI2BB2XL U1661 ( .B0(n1963), .B1(n2232), .A0N(\register[21][16] ), .A1N(
        n2233), .Y(n418) );
  OAI2BB2XL U1662 ( .B0(n1960), .B1(n2232), .A0N(\register[21][17] ), .A1N(
        n2233), .Y(n419) );
  OAI2BB2XL U1663 ( .B0(n1954), .B1(n2232), .A0N(\register[21][19] ), .A1N(
        n2233), .Y(n421) );
  OAI2BB2XL U1664 ( .B0(n1951), .B1(n2232), .A0N(\register[21][20] ), .A1N(
        n2233), .Y(n422) );
  OAI2BB2XL U1665 ( .B0(n1948), .B1(n2232), .A0N(\register[21][21] ), .A1N(
        n2232), .Y(n423) );
  OAI2BB2XL U1666 ( .B0(n1945), .B1(n2232), .A0N(\register[21][22] ), .A1N(
        n2232), .Y(n424) );
  OAI2BB2XL U1667 ( .B0(n1942), .B1(n2232), .A0N(\register[21][23] ), .A1N(
        n2232), .Y(n425) );
  OAI2BB2XL U1668 ( .B0(n1939), .B1(n2232), .A0N(\register[21][24] ), .A1N(
        n2232), .Y(n426) );
  OAI2BB2XL U1669 ( .B0(n1930), .B1(n2231), .A0N(\register[21][27] ), .A1N(
        n2232), .Y(n429) );
  OAI2BB2XL U1670 ( .B0(n1927), .B1(n2230), .A0N(\register[21][28] ), .A1N(
        n2232), .Y(n430) );
  OAI2BB2XL U1671 ( .B0(n1924), .B1(n2230), .A0N(\register[21][29] ), .A1N(
        n2232), .Y(n431) );
  OAI2BB2XL U1672 ( .B0(n1921), .B1(n2230), .A0N(\register[21][30] ), .A1N(
        n2232), .Y(n432) );
  OAI2BB2XL U1673 ( .B0(n1918), .B1(n2230), .A0N(\register[21][31] ), .A1N(
        n2232), .Y(n433) );
  OAI2BB2XL U1674 ( .B0(n2011), .B1(n2226), .A0N(\register[20][0] ), .A1N(
        n2228), .Y(n434) );
  OAI2BB2XL U1675 ( .B0(n2008), .B1(n2226), .A0N(\register[20][1] ), .A1N(
        n2229), .Y(n435) );
  OAI2BB2XL U1676 ( .B0(n2005), .B1(n2226), .A0N(\register[20][2] ), .A1N(
        n2229), .Y(n436) );
  OAI2BB2XL U1677 ( .B0(n2002), .B1(n2226), .A0N(\register[20][3] ), .A1N(
        n2229), .Y(n437) );
  OAI2BB2XL U1678 ( .B0(n1999), .B1(n2226), .A0N(\register[20][4] ), .A1N(
        n2229), .Y(n438) );
  OAI2BB2XL U1679 ( .B0(n1996), .B1(n2226), .A0N(\register[20][5] ), .A1N(
        n2229), .Y(n439) );
  OAI2BB2XL U1680 ( .B0(n1993), .B1(n2226), .A0N(\register[20][6] ), .A1N(
        n2229), .Y(n440) );
  OAI2BB2XL U1681 ( .B0(n1990), .B1(n2226), .A0N(\register[20][7] ), .A1N(
        n2229), .Y(n441) );
  OAI2BB2XL U1682 ( .B0(n1987), .B1(n2227), .A0N(\register[20][8] ), .A1N(
        n2229), .Y(n442) );
  OAI2BB2XL U1683 ( .B0(n1984), .B1(n2227), .A0N(\register[20][9] ), .A1N(
        n2229), .Y(n443) );
  OAI2BB2XL U1684 ( .B0(n1981), .B1(n2227), .A0N(\register[20][10] ), .A1N(
        n2229), .Y(n444) );
  OAI2BB2XL U1685 ( .B0(n1978), .B1(n2227), .A0N(\register[20][11] ), .A1N(
        n2229), .Y(n445) );
  OAI2BB2XL U1686 ( .B0(n1975), .B1(n2227), .A0N(\register[20][12] ), .A1N(
        n2229), .Y(n446) );
  OAI2BB2XL U1687 ( .B0(n1972), .B1(n2227), .A0N(\register[20][13] ), .A1N(
        n2229), .Y(n447) );
  OAI2BB2XL U1688 ( .B0(n1969), .B1(n2227), .A0N(\register[20][14] ), .A1N(
        n2229), .Y(n448) );
  OAI2BB2XL U1689 ( .B0(n1966), .B1(n2227), .A0N(\register[20][15] ), .A1N(
        n2229), .Y(n449) );
  OAI2BB2XL U1690 ( .B0(n1963), .B1(n2228), .A0N(\register[20][16] ), .A1N(
        n2229), .Y(n450) );
  OAI2BB2XL U1691 ( .B0(n1923), .B1(n2186), .A0N(\register[10][29] ), .A1N(
        n2188), .Y(n783) );
  OAI2BB2XL U1692 ( .B0(n1992), .B1(n2162), .A0N(\register[4][6] ), .A1N(n2165), .Y(n952) );
  OAI2BB2XL U1693 ( .B0(n1968), .B1(n2163), .A0N(\register[4][14] ), .A1N(
        n2165), .Y(n960) );
  OAI2BB2XL U1694 ( .B0(n1968), .B1(n2155), .A0N(\register[2][14] ), .A1N(
        n2157), .Y(n1024) );
  OAI2BB2XL U1695 ( .B0(n1920), .B1(n2154), .A0N(\register[2][30] ), .A1N(
        n2156), .Y(n1040) );
  OAI2BB2XL U1696 ( .B0(n1992), .B1(n2150), .A0N(\register[1][6] ), .A1N(n2153), .Y(n1048) );
  OAI2BB2XL U1697 ( .B0(n1977), .B1(n2151), .A0N(\register[1][11] ), .A1N(
        n2153), .Y(n1053) );
  OAI2BB2XL U1698 ( .B0(n1975), .B1(n2231), .A0N(\register[21][12] ), .A1N(
        n2233), .Y(n414) );
  OAI2BB2XL U1699 ( .B0(n1972), .B1(n2231), .A0N(\register[21][13] ), .A1N(
        n2233), .Y(n415) );
  OAI2BB2XL U1700 ( .B0(n1969), .B1(n2231), .A0N(\register[21][14] ), .A1N(
        n2233), .Y(n416) );
  OAI2BB2XL U1701 ( .B0(n1966), .B1(n2231), .A0N(\register[21][15] ), .A1N(
        n2233), .Y(n417) );
  OAI2BB2XL U1702 ( .B0(n1957), .B1(n2231), .A0N(\register[21][18] ), .A1N(
        n2233), .Y(n420) );
  OAI2BB2XL U1703 ( .B0(n1936), .B1(n2231), .A0N(\register[21][25] ), .A1N(
        n2232), .Y(n427) );
  OAI2BB2XL U1704 ( .B0(n1933), .B1(n2231), .A0N(\register[21][26] ), .A1N(
        n2232), .Y(n428) );
  OAI2BB2XL U1705 ( .B0(n1957), .B1(n2227), .A0N(\register[20][18] ), .A1N(
        n2229), .Y(n452) );
  OAI2BB2XL U1706 ( .B0(n1954), .B1(n2228), .A0N(\register[20][19] ), .A1N(
        n2229), .Y(n453) );
  OAI2BB2XL U1707 ( .B0(n1951), .B1(n2228), .A0N(\register[20][20] ), .A1N(
        n2229), .Y(n454) );
  OAI2BB2XL U1708 ( .B0(n1948), .B1(n2228), .A0N(\register[20][21] ), .A1N(
        n2228), .Y(n455) );
  OAI2BB2XL U1709 ( .B0(n1945), .B1(n2228), .A0N(\register[20][22] ), .A1N(
        n2228), .Y(n456) );
  OAI2BB2XL U1710 ( .B0(n1936), .B1(n2227), .A0N(\register[20][25] ), .A1N(
        n2228), .Y(n459) );
  OAI2BB2XL U1711 ( .B0(n1933), .B1(n2227), .A0N(\register[20][26] ), .A1N(
        n2228), .Y(n460) );
  OAI2BB2XL U1712 ( .B0(n1930), .B1(n2227), .A0N(\register[20][27] ), .A1N(
        n2228), .Y(n461) );
  OAI2BB2XL U1713 ( .B0(n1927), .B1(n2226), .A0N(\register[20][28] ), .A1N(
        n2228), .Y(n462) );
  OAI2BB2XL U1714 ( .B0(n1924), .B1(n2226), .A0N(\register[20][29] ), .A1N(
        n2228), .Y(n463) );
  OAI2BB2XL U1715 ( .B0(n1921), .B1(n2226), .A0N(\register[20][30] ), .A1N(
        n2228), .Y(n464) );
  OAI2BB2XL U1716 ( .B0(n1918), .B1(n2226), .A0N(\register[20][31] ), .A1N(
        n2228), .Y(n465) );
  OAI2BB2XL U1717 ( .B0(n2011), .B1(n2222), .A0N(\register[19][0] ), .A1N(
        n2224), .Y(n466) );
  OAI2BB2XL U1718 ( .B0(n2008), .B1(n2222), .A0N(\register[19][1] ), .A1N(
        n2225), .Y(n467) );
  OAI2BB2XL U1719 ( .B0(n2005), .B1(n2222), .A0N(\register[19][2] ), .A1N(
        n2225), .Y(n468) );
  OAI2BB2XL U1720 ( .B0(n2002), .B1(n2222), .A0N(\register[19][3] ), .A1N(
        n2225), .Y(n469) );
  OAI2BB2XL U1721 ( .B0(n1999), .B1(n2222), .A0N(\register[19][4] ), .A1N(
        n2225), .Y(n470) );
  OAI2BB2XL U1722 ( .B0(n1996), .B1(n2222), .A0N(\register[19][5] ), .A1N(
        n2225), .Y(n471) );
  OAI2BB2XL U1723 ( .B0(n1993), .B1(n2222), .A0N(\register[19][6] ), .A1N(
        n2225), .Y(n472) );
  OAI2BB2XL U1724 ( .B0(n1990), .B1(n2222), .A0N(\register[19][7] ), .A1N(
        n2225), .Y(n473) );
  OAI2BB2XL U1725 ( .B0(n1987), .B1(n2223), .A0N(\register[19][8] ), .A1N(
        n2225), .Y(n474) );
  OAI2BB2XL U1726 ( .B0(n1984), .B1(n2223), .A0N(\register[19][9] ), .A1N(
        n2225), .Y(n475) );
  OAI2BB2XL U1727 ( .B0(n1981), .B1(n2223), .A0N(\register[19][10] ), .A1N(
        n2225), .Y(n476) );
  OAI2BB2XL U1728 ( .B0(n1978), .B1(n2223), .A0N(\register[19][11] ), .A1N(
        n2225), .Y(n477) );
  OAI2BB2XL U1729 ( .B0(n1975), .B1(n2223), .A0N(\register[19][12] ), .A1N(
        n2225), .Y(n478) );
  OAI2BB2XL U1730 ( .B0(n1972), .B1(n2223), .A0N(\register[19][13] ), .A1N(
        n2225), .Y(n479) );
  OAI2BB2XL U1731 ( .B0(n1969), .B1(n2223), .A0N(\register[19][14] ), .A1N(
        n2225), .Y(n480) );
  OAI2BB2XL U1732 ( .B0(n1966), .B1(n2223), .A0N(\register[19][15] ), .A1N(
        n2225), .Y(n481) );
  OAI2BB2XL U1733 ( .B0(n1963), .B1(n2224), .A0N(\register[19][16] ), .A1N(
        n2225), .Y(n482) );
  OAI2BB2XL U1734 ( .B0(n1960), .B1(n2224), .A0N(\register[19][17] ), .A1N(
        n2225), .Y(n483) );
  OAI2BB2XL U1735 ( .B0(n1951), .B1(n2224), .A0N(\register[19][20] ), .A1N(
        n2225), .Y(n486) );
  OAI2BB2XL U1736 ( .B0(n1948), .B1(n2224), .A0N(\register[19][21] ), .A1N(
        n2224), .Y(n487) );
  OAI2BB2XL U1737 ( .B0(n1945), .B1(n2224), .A0N(\register[19][22] ), .A1N(
        n2224), .Y(n488) );
  OAI2BB2XL U1738 ( .B0(n1942), .B1(n2224), .A0N(\register[19][23] ), .A1N(
        n2224), .Y(n489) );
  OAI2BB2XL U1739 ( .B0(n1939), .B1(n2224), .A0N(\register[19][24] ), .A1N(
        n2224), .Y(n490) );
  OAI2BB2XL U1740 ( .B0(n2004), .B1(n2182), .A0N(\register[9][2] ), .A1N(n2185), .Y(n788) );
  OAI2BB2XL U1741 ( .B0(n2001), .B1(n2182), .A0N(\register[9][3] ), .A1N(n2185), .Y(n789) );
  OAI2BB2XL U1742 ( .B0(n1962), .B1(n2184), .A0N(\register[9][16] ), .A1N(
        n2185), .Y(n802) );
  OAI2BB2XL U1743 ( .B0(n1956), .B1(n2183), .A0N(\register[9][18] ), .A1N(
        n2185), .Y(n804) );
  OAI2BB2XL U1744 ( .B0(n1929), .B1(n2183), .A0N(\register[9][27] ), .A1N(
        n2184), .Y(n813) );
  OAI2BB2XL U1745 ( .B0(n1917), .B1(n2182), .A0N(\register[9][31] ), .A1N(
        n2184), .Y(n817) );
  OAI2BB2XL U1746 ( .B0(n1923), .B1(n2162), .A0N(\register[4][29] ), .A1N(
        n2164), .Y(n975) );
  OAI2BB2XL U1747 ( .B0(n2004), .B1(n2158), .A0N(\register[3][2] ), .A1N(n2161), .Y(n980) );
  OAI2BB2XL U1748 ( .B0(n1962), .B1(n2152), .A0N(\register[1][16] ), .A1N(
        n2153), .Y(n1058) );
  OAI2BB2XL U1749 ( .B0(n1942), .B1(n2228), .A0N(\register[20][23] ), .A1N(
        n2228), .Y(n457) );
  OAI2BB2XL U1750 ( .B0(n1932), .B1(n2163), .A0N(\register[4][26] ), .A1N(
        n2164), .Y(n972) );
  OAI2BB2XL U1751 ( .B0(n1965), .B1(n2151), .A0N(\register[1][15] ), .A1N(
        n2153), .Y(n1057) );
  OAI2BB2XL U1752 ( .B0(n1932), .B1(n2147), .A0N(\register[0][26] ), .A1N(
        n2148), .Y(n1100) );
  OAI2BB2XL U1753 ( .B0(n1929), .B1(n2147), .A0N(\register[0][27] ), .A1N(
        n2148), .Y(n1101) );
  OAI2BB2XL U1754 ( .B0(n1957), .B1(n2223), .A0N(\register[19][18] ), .A1N(
        n2225), .Y(n484) );
  OAI2BB2XL U1755 ( .B0(n1936), .B1(n2223), .A0N(\register[19][25] ), .A1N(
        n2224), .Y(n491) );
  OAI2BB2XL U1756 ( .B0(n1933), .B1(n2223), .A0N(\register[19][26] ), .A1N(
        n2224), .Y(n492) );
  OAI2BB2XL U1757 ( .B0(n1930), .B1(n2223), .A0N(\register[19][27] ), .A1N(
        n2224), .Y(n493) );
  OAI2BB2XL U1758 ( .B0(n1927), .B1(n2222), .A0N(\register[19][28] ), .A1N(
        n2224), .Y(n494) );
  OAI2BB2XL U1759 ( .B0(n1924), .B1(n2222), .A0N(\register[19][29] ), .A1N(
        n2224), .Y(n495) );
  OAI2BB2XL U1760 ( .B0(n1921), .B1(n2222), .A0N(\register[19][30] ), .A1N(
        n2224), .Y(n496) );
  OAI2BB2XL U1761 ( .B0(n1918), .B1(n2222), .A0N(\register[19][31] ), .A1N(
        n2224), .Y(n497) );
  OAI2BB2XL U1762 ( .B0(n2011), .B1(n2218), .A0N(\register[18][0] ), .A1N(
        n2220), .Y(n498) );
  OAI2BB2XL U1763 ( .B0(n2008), .B1(n2218), .A0N(\register[18][1] ), .A1N(
        n2221), .Y(n499) );
  OAI2BB2XL U1764 ( .B0(n2005), .B1(n2218), .A0N(\register[18][2] ), .A1N(
        n2221), .Y(n500) );
  OAI2BB2XL U1765 ( .B0(n2002), .B1(n2218), .A0N(\register[18][3] ), .A1N(
        n2221), .Y(n501) );
  OAI2BB2XL U1766 ( .B0(n1999), .B1(n2218), .A0N(\register[18][4] ), .A1N(
        n2221), .Y(n502) );
  OAI2BB2XL U1767 ( .B0(n1963), .B1(n2220), .A0N(\register[18][16] ), .A1N(
        n2221), .Y(n514) );
  OAI2BB2XL U1768 ( .B0(n1960), .B1(n2220), .A0N(\register[18][17] ), .A1N(
        n2221), .Y(n515) );
  OAI2BB2XL U1769 ( .B0(n1935), .B1(n2151), .A0N(\register[1][25] ), .A1N(
        n2152), .Y(n1067) );
  OAI2BB2XL U1770 ( .B0(n1917), .B1(n2146), .A0N(\register[0][31] ), .A1N(
        n2148), .Y(n1105) );
  OAI2BB2XL U1771 ( .B0(n1996), .B1(n2218), .A0N(\register[18][5] ), .A1N(
        n2221), .Y(n503) );
  OAI2BB2XL U1772 ( .B0(n1993), .B1(n2218), .A0N(\register[18][6] ), .A1N(
        n2221), .Y(n504) );
  OAI2BB2XL U1773 ( .B0(n1990), .B1(n2218), .A0N(\register[18][7] ), .A1N(
        n2221), .Y(n505) );
  OAI2BB2XL U1774 ( .B0(n1987), .B1(n2219), .A0N(\register[18][8] ), .A1N(
        n2221), .Y(n506) );
  OAI2BB2XL U1775 ( .B0(n1984), .B1(n2219), .A0N(\register[18][9] ), .A1N(
        n2221), .Y(n507) );
  OAI2BB2XL U1776 ( .B0(n1981), .B1(n2219), .A0N(\register[18][10] ), .A1N(
        n2221), .Y(n508) );
  OAI2BB2XL U1777 ( .B0(n1978), .B1(n2219), .A0N(\register[18][11] ), .A1N(
        n2221), .Y(n509) );
  OAI2BB2XL U1778 ( .B0(n1975), .B1(n2219), .A0N(\register[18][12] ), .A1N(
        n2221), .Y(n510) );
  OAI2BB2XL U1779 ( .B0(n1972), .B1(n2219), .A0N(\register[18][13] ), .A1N(
        n2221), .Y(n511) );
  OAI2BB2XL U1780 ( .B0(n1969), .B1(n2219), .A0N(\register[18][14] ), .A1N(
        n2221), .Y(n512) );
  OAI2BB2XL U1781 ( .B0(n1966), .B1(n2219), .A0N(\register[18][15] ), .A1N(
        n2221), .Y(n513) );
  OAI2BB2XL U1782 ( .B0(n1957), .B1(n2219), .A0N(\register[18][18] ), .A1N(
        n2221), .Y(n516) );
  OAI2BB2XL U1783 ( .B0(n1936), .B1(n2219), .A0N(\register[18][25] ), .A1N(
        n2220), .Y(n523) );
  OAI2BB2XL U1784 ( .B0(n1933), .B1(n2219), .A0N(\register[18][26] ), .A1N(
        n2220), .Y(n524) );
  OAI2BB2XL U1785 ( .B0(n1930), .B1(n2219), .A0N(\register[18][27] ), .A1N(
        n2220), .Y(n525) );
  OAI2BB2XL U1786 ( .B0(n1927), .B1(n2218), .A0N(\register[18][28] ), .A1N(
        n2220), .Y(n526) );
  OAI2BB2XL U1787 ( .B0(n1924), .B1(n2218), .A0N(\register[18][29] ), .A1N(
        n2220), .Y(n527) );
  OAI2BB2XL U1788 ( .B0(n1921), .B1(n2218), .A0N(\register[18][30] ), .A1N(
        n2220), .Y(n528) );
  OAI2BB2XL U1789 ( .B0(n1918), .B1(n2218), .A0N(\register[18][31] ), .A1N(
        n2220), .Y(n529) );
  OAI2BB2XL U1790 ( .B0(n2011), .B1(n2214), .A0N(\register[17][0] ), .A1N(
        n2216), .Y(n530) );
  OAI2BB2XL U1791 ( .B0(n2008), .B1(n2214), .A0N(\register[17][1] ), .A1N(
        n2217), .Y(n531) );
  OAI2BB2XL U1792 ( .B0(n2005), .B1(n2214), .A0N(\register[17][2] ), .A1N(
        n2217), .Y(n532) );
  OAI2BB2XL U1793 ( .B0(n2002), .B1(n2214), .A0N(\register[17][3] ), .A1N(
        n2217), .Y(n533) );
  OAI2BB2XL U1794 ( .B0(n1999), .B1(n2214), .A0N(\register[17][4] ), .A1N(
        n2217), .Y(n534) );
  OAI2BB2XL U1795 ( .B0(n1996), .B1(n2214), .A0N(\register[17][5] ), .A1N(
        n2217), .Y(n535) );
  OAI2BB2XL U1796 ( .B0(n1993), .B1(n2214), .A0N(\register[17][6] ), .A1N(
        n2217), .Y(n536) );
  OAI2BB2XL U1797 ( .B0(n1990), .B1(n2214), .A0N(\register[17][7] ), .A1N(
        n2217), .Y(n537) );
  OAI2BB2XL U1798 ( .B0(n1987), .B1(n2215), .A0N(\register[17][8] ), .A1N(
        n2217), .Y(n538) );
  OAI2BB2XL U1799 ( .B0(n1984), .B1(n2215), .A0N(\register[17][9] ), .A1N(
        n2217), .Y(n539) );
  OAI2BB2XL U1800 ( .B0(n1963), .B1(n2216), .A0N(\register[17][16] ), .A1N(
        n2217), .Y(n546) );
  OAI2BB2XL U1801 ( .B0(n1960), .B1(n2216), .A0N(\register[17][17] ), .A1N(
        n2217), .Y(n547) );
  OAI2BB2XL U1802 ( .B0(n2001), .B1(n2158), .A0N(\register[3][3] ), .A1N(n2161), .Y(n981) );
  OAI2BB2XL U1803 ( .B0(n1974), .B1(n2159), .A0N(\register[3][12] ), .A1N(
        n2161), .Y(n990) );
  OAI2BB2XL U1804 ( .B0(n1971), .B1(n2151), .A0N(\register[1][13] ), .A1N(
        n2153), .Y(n1055) );
  OAI2BB2XL U1805 ( .B0(n1932), .B1(n2151), .A0N(\register[1][26] ), .A1N(
        n2152), .Y(n1068) );
  OAI2BB2XL U1806 ( .B0(n1920), .B1(n2146), .A0N(\register[0][30] ), .A1N(
        n2148), .Y(n1104) );
  OAI2BB2XL U1807 ( .B0(n1981), .B1(n2215), .A0N(\register[17][10] ), .A1N(
        n2217), .Y(n540) );
  OAI2BB2XL U1808 ( .B0(n1978), .B1(n2215), .A0N(\register[17][11] ), .A1N(
        n2217), .Y(n541) );
  OAI2BB2XL U1809 ( .B0(n1975), .B1(n2215), .A0N(\register[17][12] ), .A1N(
        n2217), .Y(n542) );
  OAI2BB2XL U1810 ( .B0(n1972), .B1(n2215), .A0N(\register[17][13] ), .A1N(
        n2217), .Y(n543) );
  OAI2BB2XL U1811 ( .B0(n1969), .B1(n2215), .A0N(\register[17][14] ), .A1N(
        n2217), .Y(n544) );
  OAI2BB2XL U1812 ( .B0(n1966), .B1(n2215), .A0N(\register[17][15] ), .A1N(
        n2217), .Y(n545) );
  OAI2BB2XL U1813 ( .B0(n1957), .B1(n2215), .A0N(\register[17][18] ), .A1N(
        n2217), .Y(n548) );
  OAI2BB2XL U1814 ( .B0(n1954), .B1(n2216), .A0N(\register[17][19] ), .A1N(
        n2217), .Y(n549) );
  OAI2BB2XL U1815 ( .B0(n1951), .B1(n2216), .A0N(\register[17][20] ), .A1N(
        n2217), .Y(n550) );
  OAI2BB2XL U1816 ( .B0(n1948), .B1(n2216), .A0N(\register[17][21] ), .A1N(
        n2216), .Y(n551) );
  OAI2BB2XL U1817 ( .B0(n1945), .B1(n2216), .A0N(\register[17][22] ), .A1N(
        n2216), .Y(n552) );
  OAI2BB2XL U1818 ( .B0(n1942), .B1(n2216), .A0N(\register[17][23] ), .A1N(
        n2216), .Y(n553) );
  OAI2BB2XL U1819 ( .B0(n1939), .B1(n2216), .A0N(\register[17][24] ), .A1N(
        n2216), .Y(n554) );
  OAI2BB2XL U1820 ( .B0(n1936), .B1(n2215), .A0N(\register[17][25] ), .A1N(
        n2216), .Y(n555) );
  OAI2BB2XL U1821 ( .B0(n1933), .B1(n2215), .A0N(\register[17][26] ), .A1N(
        n2216), .Y(n556) );
  OAI2BB2XL U1822 ( .B0(n1930), .B1(n2215), .A0N(\register[17][27] ), .A1N(
        n2216), .Y(n557) );
  OAI2BB2XL U1823 ( .B0(n1927), .B1(n2214), .A0N(\register[17][28] ), .A1N(
        n2216), .Y(n558) );
  OAI2BB2XL U1824 ( .B0(n1924), .B1(n2214), .A0N(\register[17][29] ), .A1N(
        n2216), .Y(n559) );
  OAI2BB2XL U1825 ( .B0(n1921), .B1(n2214), .A0N(\register[17][30] ), .A1N(
        n2216), .Y(n560) );
  OAI2BB2XL U1826 ( .B0(n1918), .B1(n2214), .A0N(\register[17][31] ), .A1N(
        n2216), .Y(n561) );
  OAI2BB2XL U1827 ( .B0(n2011), .B1(n2210), .A0N(\register[16][0] ), .A1N(
        n2212), .Y(n562) );
  OAI2BB2XL U1828 ( .B0(n2008), .B1(n2210), .A0N(\register[16][1] ), .A1N(
        n2213), .Y(n563) );
  OAI2BB2XL U1829 ( .B0(n2005), .B1(n2210), .A0N(\register[16][2] ), .A1N(
        n2213), .Y(n564) );
  OAI2BB2XL U1830 ( .B0(n2002), .B1(n2210), .A0N(\register[16][3] ), .A1N(
        n2213), .Y(n565) );
  OAI2BB2XL U1831 ( .B0(n1999), .B1(n2210), .A0N(\register[16][4] ), .A1N(
        n2213), .Y(n566) );
  OAI2BB2XL U1832 ( .B0(n1996), .B1(n2210), .A0N(\register[16][5] ), .A1N(
        n2213), .Y(n567) );
  OAI2BB2XL U1833 ( .B0(n1993), .B1(n2210), .A0N(\register[16][6] ), .A1N(
        n2213), .Y(n568) );
  OAI2BB2XL U1834 ( .B0(n1990), .B1(n2210), .A0N(\register[16][7] ), .A1N(
        n2213), .Y(n569) );
  OAI2BB2XL U1835 ( .B0(n1987), .B1(n2211), .A0N(\register[16][8] ), .A1N(
        n2213), .Y(n570) );
  OAI2BB2XL U1836 ( .B0(n1984), .B1(n2211), .A0N(\register[16][9] ), .A1N(
        n2213), .Y(n571) );
  OAI2BB2XL U1837 ( .B0(n1981), .B1(n2211), .A0N(\register[16][10] ), .A1N(
        n2213), .Y(n572) );
  OAI2BB2XL U1838 ( .B0(n1978), .B1(n2211), .A0N(\register[16][11] ), .A1N(
        n2213), .Y(n573) );
  OAI2BB2XL U1839 ( .B0(n1975), .B1(n2211), .A0N(\register[16][12] ), .A1N(
        n2213), .Y(n574) );
  OAI2BB2XL U1840 ( .B0(n1972), .B1(n2211), .A0N(\register[16][13] ), .A1N(
        n2213), .Y(n575) );
  OAI2BB2XL U1841 ( .B0(n1969), .B1(n2211), .A0N(\register[16][14] ), .A1N(
        n2213), .Y(n576) );
  OAI2BB2XL U1842 ( .B0(n1966), .B1(n2211), .A0N(\register[16][15] ), .A1N(
        n2213), .Y(n577) );
  OAI2BB2XL U1843 ( .B0(n1957), .B1(n2211), .A0N(\register[16][18] ), .A1N(
        n2213), .Y(n580) );
  OAI2BB2XL U1844 ( .B0(n1936), .B1(n2211), .A0N(\register[16][25] ), .A1N(
        n2212), .Y(n587) );
  OAI2BB2XL U1845 ( .B0(n1933), .B1(n2211), .A0N(\register[16][26] ), .A1N(
        n2212), .Y(n588) );
  OAI2BB2XL U1846 ( .B0(n1930), .B1(n2211), .A0N(\register[16][27] ), .A1N(
        n2212), .Y(n589) );
  OAI2BB2XL U1847 ( .B0(n1927), .B1(n2210), .A0N(\register[16][28] ), .A1N(
        n2212), .Y(n590) );
  OAI2BB2XL U1848 ( .B0(n1924), .B1(n2210), .A0N(\register[16][29] ), .A1N(
        n2212), .Y(n591) );
  OAI2BB2XL U1849 ( .B0(n1921), .B1(n2210), .A0N(\register[16][30] ), .A1N(
        n2212), .Y(n592) );
  OAI2BB2XL U1850 ( .B0(n1918), .B1(n2210), .A0N(\register[16][31] ), .A1N(
        n2212), .Y(n593) );
  OAI2BB2XL U1851 ( .B0(n2270), .B1(n2012), .A0N(\register[31][0] ), .A1N(
        n2272), .Y(n82) );
  OAI2BB2XL U1852 ( .B0(n2270), .B1(n2009), .A0N(\register[31][1] ), .A1N(
        n2273), .Y(n83) );
  OAI2BB2XL U1853 ( .B0(n2270), .B1(n2006), .A0N(\register[31][2] ), .A1N(
        n2273), .Y(n84) );
  OAI2BB2XL U1854 ( .B0(n2270), .B1(n2003), .A0N(\register[31][3] ), .A1N(
        n2273), .Y(n85) );
  OAI2BB2XL U1855 ( .B0(n2270), .B1(n2000), .A0N(\register[31][4] ), .A1N(
        n2273), .Y(n86) );
  OAI2BB2XL U1856 ( .B0(n2270), .B1(n1997), .A0N(\register[31][5] ), .A1N(
        n2273), .Y(n87) );
  OAI2BB2XL U1857 ( .B0(n2270), .B1(n1994), .A0N(\register[31][6] ), .A1N(
        n2273), .Y(n88) );
  OAI2BB2XL U1858 ( .B0(n2270), .B1(n1991), .A0N(\register[31][7] ), .A1N(
        n2273), .Y(n89) );
  OAI2BB2XL U1859 ( .B0(n2271), .B1(n1988), .A0N(\register[31][8] ), .A1N(
        n2273), .Y(n90) );
  OAI2BB2XL U1860 ( .B0(n2271), .B1(n1985), .A0N(\register[31][9] ), .A1N(
        n2273), .Y(n91) );
  OAI2BB2XL U1861 ( .B0(n2271), .B1(n1982), .A0N(\register[31][10] ), .A1N(
        n2273), .Y(n92) );
  OAI2BB2XL U1862 ( .B0(n2271), .B1(n1979), .A0N(\register[31][11] ), .A1N(
        n2273), .Y(n93) );
  OAI2BB2XL U1863 ( .B0(n2271), .B1(n1976), .A0N(\register[31][12] ), .A1N(
        n2273), .Y(n94) );
  OAI2BB2XL U1864 ( .B0(n2271), .B1(n1973), .A0N(\register[31][13] ), .A1N(
        n2273), .Y(n95) );
  OAI2BB2XL U1865 ( .B0(n2271), .B1(n1970), .A0N(\register[31][14] ), .A1N(
        n2273), .Y(n96) );
  OAI2BB2XL U1866 ( .B0(n2271), .B1(n1967), .A0N(\register[31][15] ), .A1N(
        n2273), .Y(n97) );
  OAI2BB2XL U1867 ( .B0(n2272), .B1(n1964), .A0N(\register[31][16] ), .A1N(
        n2273), .Y(n98) );
  OAI2BB2XL U1868 ( .B0(n2272), .B1(n1961), .A0N(\register[31][17] ), .A1N(
        n2273), .Y(n99) );
  OAI2BB2XL U1869 ( .B0(n2271), .B1(n1958), .A0N(\register[31][18] ), .A1N(
        n2273), .Y(n100) );
  OAI2BB2XL U1870 ( .B0(n2272), .B1(n1955), .A0N(\register[31][19] ), .A1N(
        n2273), .Y(n101) );
  OAI2BB2XL U1871 ( .B0(n2272), .B1(n1952), .A0N(\register[31][20] ), .A1N(
        n2272), .Y(n102) );
  OAI2BB2XL U1872 ( .B0(n2272), .B1(n1949), .A0N(\register[31][21] ), .A1N(
        n2272), .Y(n103) );
  OAI2BB2XL U1873 ( .B0(n2272), .B1(n1946), .A0N(\register[31][22] ), .A1N(
        n2272), .Y(n104) );
  OAI2BB2XL U1874 ( .B0(n2272), .B1(n1943), .A0N(\register[31][23] ), .A1N(
        n2272), .Y(n105) );
  OAI2BB2XL U1875 ( .B0(n2272), .B1(n1940), .A0N(\register[31][24] ), .A1N(
        n2272), .Y(n106) );
  OAI2BB2XL U1876 ( .B0(n2271), .B1(n1937), .A0N(\register[31][25] ), .A1N(
        n2272), .Y(n107) );
  OAI2BB2XL U1877 ( .B0(n2271), .B1(n1934), .A0N(\register[31][26] ), .A1N(
        n2272), .Y(n108) );
  OAI2BB2XL U1878 ( .B0(n2271), .B1(n1931), .A0N(\register[31][27] ), .A1N(
        n2272), .Y(n109) );
  OAI2BB2XL U1879 ( .B0(n2270), .B1(n1928), .A0N(\register[31][28] ), .A1N(
        n2272), .Y(n110) );
  OAI2BB2XL U1880 ( .B0(n2270), .B1(n1925), .A0N(\register[31][29] ), .A1N(
        n2272), .Y(n111) );
  OAI2BB2XL U1881 ( .B0(n2270), .B1(n1922), .A0N(\register[31][30] ), .A1N(
        n2272), .Y(n112) );
  OAI2BB2XL U1882 ( .B0(n2270), .B1(n1919), .A0N(\register[31][31] ), .A1N(
        n2272), .Y(n113) );
  MXI2X1 U1883 ( .A(n1511), .B(n1512), .S0(n1814), .Y(ReadData2_o[9]) );
  MX4X1 U1884 ( .A(n1632), .B(n1630), .C(n1631), .D(n1629), .S0(n1820), .S1(
        n1828), .Y(n1512) );
  MX4X1 U1885 ( .A(n1636), .B(n1634), .C(n1635), .D(n1633), .S0(n1820), .S1(
        n1828), .Y(n1511) );
  MXI4X1 U1886 ( .A(\register[28][9] ), .B(\register[29][9] ), .C(
        \register[30][9] ), .D(\register[31][9] ), .S0(n1899), .S1(n1858), .Y(
        n1629) );
  MXI2X1 U1887 ( .A(n1513), .B(n1514), .S0(n1814), .Y(ReadData2_o[10]) );
  MX4X1 U1888 ( .A(n1640), .B(n1638), .C(n1639), .D(n1637), .S0(n1820), .S1(
        n1828), .Y(n1514) );
  MX4X1 U1889 ( .A(n1644), .B(n1642), .C(n1643), .D(n1641), .S0(n1820), .S1(
        n1828), .Y(n1513) );
  MXI4X1 U1890 ( .A(\register[28][10] ), .B(\register[29][10] ), .C(
        \register[30][10] ), .D(\register[31][10] ), .S0(n1900), .S1(n1859), 
        .Y(n1637) );
  MXI2X1 U1891 ( .A(n1515), .B(n1516), .S0(n1814), .Y(ReadData2_o[11]) );
  MX4X1 U1892 ( .A(n1648), .B(n1646), .C(n1647), .D(n1645), .S0(n1820), .S1(
        n1828), .Y(n1516) );
  MX4X1 U1893 ( .A(n1652), .B(n1650), .C(n1651), .D(n1649), .S0(n1820), .S1(
        n1828), .Y(n1515) );
  MXI4X1 U1894 ( .A(\register[28][11] ), .B(\register[29][11] ), .C(
        \register[30][11] ), .D(\register[31][11] ), .S0(n1901), .S1(n1860), 
        .Y(n1645) );
  MXI2X1 U1895 ( .A(n1517), .B(n1518), .S0(n1814), .Y(ReadData2_o[12]) );
  MX4X1 U1896 ( .A(n1656), .B(n1654), .C(n1655), .D(n1653), .S0(n1820), .S1(
        n1828), .Y(n1518) );
  MX4X1 U1897 ( .A(n1660), .B(n1658), .C(n1659), .D(n1657), .S0(n1820), .S1(
        n1829), .Y(n1517) );
  MXI4X1 U1898 ( .A(\register[28][12] ), .B(\register[29][12] ), .C(
        \register[30][12] ), .D(\register[31][12] ), .S0(n1901), .S1(n1860), 
        .Y(n1653) );
  MXI2X1 U1899 ( .A(n1519), .B(n1520), .S0(n1814), .Y(ReadData2_o[13]) );
  MX4X1 U1900 ( .A(n1664), .B(n1662), .C(n1663), .D(n1661), .S0(n1820), .S1(
        n1829), .Y(n1520) );
  MX4X1 U1901 ( .A(n1668), .B(n1666), .C(n1667), .D(n1665), .S0(n1820), .S1(
        n1829), .Y(n1519) );
  MXI4X1 U1902 ( .A(\register[28][13] ), .B(\register[29][13] ), .C(
        \register[30][13] ), .D(\register[31][13] ), .S0(n1902), .S1(n1861), 
        .Y(n1661) );
  MXI2X1 U1903 ( .A(n1521), .B(n1522), .S0(n1814), .Y(ReadData2_o[14]) );
  MX4X1 U1904 ( .A(n1672), .B(n1670), .C(n1671), .D(n1669), .S0(n1821), .S1(
        n1829), .Y(n1522) );
  MX4X1 U1905 ( .A(n1676), .B(n1674), .C(n1675), .D(n1673), .S0(n1821), .S1(
        n1829), .Y(n1521) );
  MXI4X1 U1906 ( .A(\register[28][14] ), .B(\register[29][14] ), .C(
        \register[30][14] ), .D(\register[31][14] ), .S0(n1903), .S1(n1862), 
        .Y(n1669) );
  MXI2X1 U1907 ( .A(n1523), .B(n1524), .S0(n1814), .Y(ReadData2_o[15]) );
  MX4X1 U1908 ( .A(n1680), .B(n1678), .C(n1679), .D(n1677), .S0(n1821), .S1(
        n1829), .Y(n1524) );
  MX4X1 U1909 ( .A(n1684), .B(n1682), .C(n1683), .D(n1681), .S0(n1821), .S1(
        n1829), .Y(n1523) );
  MXI4X1 U1910 ( .A(\register[28][15] ), .B(\register[29][15] ), .C(
        \register[30][15] ), .D(\register[31][15] ), .S0(n1903), .S1(n1862), 
        .Y(n1677) );
  MXI2X1 U1911 ( .A(n1525), .B(n1526), .S0(n1814), .Y(ReadData2_o[16]) );
  MX4X1 U1912 ( .A(n1688), .B(n1686), .C(n1687), .D(n1685), .S0(n1821), .S1(
        n1829), .Y(n1526) );
  MX4X1 U1913 ( .A(n1692), .B(n1690), .C(n1691), .D(n1689), .S0(n1821), .S1(
        n1829), .Y(n1525) );
  MXI4X1 U1914 ( .A(\register[28][16] ), .B(\register[29][16] ), .C(
        \register[30][16] ), .D(\register[31][16] ), .S0(n1904), .S1(n1863), 
        .Y(n1685) );
  MXI2X1 U1915 ( .A(n1527), .B(n1528), .S0(n1814), .Y(ReadData2_o[17]) );
  MX4X1 U1916 ( .A(n1696), .B(n1694), .C(n1695), .D(n1693), .S0(n1821), .S1(
        n1829), .Y(n1528) );
  MX4X1 U1917 ( .A(n1700), .B(n1698), .C(n1699), .D(n1697), .S0(n1821), .S1(
        n1829), .Y(n1527) );
  MXI4X1 U1918 ( .A(\register[28][17] ), .B(\register[29][17] ), .C(
        \register[30][17] ), .D(\register[31][17] ), .S0(n1905), .S1(n1864), 
        .Y(n1693) );
  MXI2X1 U1919 ( .A(n1529), .B(n1530), .S0(n1814), .Y(ReadData2_o[18]) );
  MX4X1 U1920 ( .A(n1704), .B(n1702), .C(n1703), .D(n1701), .S0(n1821), .S1(
        n1829), .Y(n1530) );
  MX4X1 U1921 ( .A(n1708), .B(n1706), .C(n1707), .D(n1705), .S0(n1821), .S1(
        n1829), .Y(n1529) );
  MXI4X1 U1922 ( .A(\register[28][18] ), .B(\register[29][18] ), .C(
        \register[30][18] ), .D(\register[31][18] ), .S0(n1905), .S1(n1864), 
        .Y(n1701) );
  MXI2X1 U1923 ( .A(n1531), .B(n1532), .S0(n1814), .Y(ReadData2_o[19]) );
  MX4X1 U1924 ( .A(n1712), .B(n1710), .C(n1711), .D(n1709), .S0(n1821), .S1(
        n1830), .Y(n1532) );
  MX4X1 U1925 ( .A(n1716), .B(n1714), .C(n1715), .D(n1713), .S0(n1821), .S1(
        n1830), .Y(n1531) );
  MXI4X1 U1926 ( .A(\register[28][19] ), .B(\register[29][19] ), .C(
        \register[30][19] ), .D(\register[31][19] ), .S0(n1906), .S1(n1865), 
        .Y(n1709) );
  MXI2X1 U1927 ( .A(n1533), .B(n1534), .S0(n1815), .Y(ReadData2_o[20]) );
  MX4X1 U1928 ( .A(n1720), .B(n1718), .C(n1719), .D(n1717), .S0(n1822), .S1(
        n1830), .Y(n1534) );
  MX4X1 U1929 ( .A(n1724), .B(n1722), .C(n1723), .D(n1721), .S0(n1822), .S1(
        n1830), .Y(n1533) );
  MXI4X1 U1930 ( .A(\register[28][20] ), .B(\register[29][20] ), .C(
        \register[30][20] ), .D(\register[31][20] ), .S0(n1907), .S1(n1866), 
        .Y(n1717) );
  MXI2X1 U1931 ( .A(n1535), .B(n1536), .S0(n1815), .Y(ReadData2_o[21]) );
  MX4X1 U1932 ( .A(n1728), .B(n1726), .C(n1727), .D(n1725), .S0(n1822), .S1(
        n1830), .Y(n1536) );
  MX4X1 U1933 ( .A(n1732), .B(n1730), .C(n1731), .D(n1729), .S0(n1822), .S1(
        n1830), .Y(n1535) );
  MXI4X1 U1934 ( .A(\register[28][21] ), .B(\register[29][21] ), .C(
        \register[30][21] ), .D(\register[31][21] ), .S0(n1907), .S1(n1866), 
        .Y(n1725) );
  MXI2X1 U1935 ( .A(n1537), .B(n1538), .S0(n1815), .Y(ReadData2_o[22]) );
  MX4X1 U1936 ( .A(n1736), .B(n1734), .C(n1735), .D(n1733), .S0(n1822), .S1(
        n1830), .Y(n1538) );
  MX4X1 U1937 ( .A(n1740), .B(n1738), .C(n1739), .D(n1737), .S0(n1822), .S1(
        n1830), .Y(n1537) );
  MXI4X1 U1938 ( .A(\register[28][22] ), .B(\register[29][22] ), .C(
        \register[30][22] ), .D(\register[31][22] ), .S0(n1908), .S1(n1867), 
        .Y(n1733) );
  MXI2X1 U1939 ( .A(n1539), .B(n1540), .S0(n1815), .Y(ReadData2_o[23]) );
  MX4X1 U1940 ( .A(n1744), .B(n1742), .C(n1743), .D(n1741), .S0(n1822), .S1(
        n1830), .Y(n1540) );
  MX4X1 U1941 ( .A(n1748), .B(n1746), .C(n1747), .D(n1745), .S0(n1822), .S1(
        n1830), .Y(n1539) );
  MXI4X1 U1942 ( .A(\register[28][23] ), .B(\register[29][23] ), .C(
        \register[30][23] ), .D(\register[31][23] ), .S0(n1909), .S1(n1868), 
        .Y(n1741) );
  MXI2X1 U1943 ( .A(n1541), .B(n1542), .S0(n1815), .Y(ReadData2_o[24]) );
  MX4X1 U1944 ( .A(n1752), .B(n1750), .C(n1751), .D(n1749), .S0(n1822), .S1(
        n1830), .Y(n1542) );
  MX4X1 U1945 ( .A(n1756), .B(n1754), .C(n1755), .D(n1753), .S0(n1822), .S1(
        n1830), .Y(n1541) );
  MXI4X1 U1946 ( .A(\register[28][24] ), .B(\register[29][24] ), .C(
        \register[30][24] ), .D(\register[31][24] ), .S0(n1909), .S1(n1868), 
        .Y(n1749) );
  MXI2X1 U1947 ( .A(n1543), .B(n1544), .S0(n1815), .Y(ReadData2_o[25]) );
  MX4X1 U1948 ( .A(n1760), .B(n1758), .C(n1759), .D(n1757), .S0(n1822), .S1(
        n1830), .Y(n1544) );
  MX4X1 U1949 ( .A(n1764), .B(n1762), .C(n1763), .D(n1761), .S0(n1822), .S1(
        n1831), .Y(n1543) );
  MXI4X1 U1950 ( .A(\register[28][25] ), .B(\register[29][25] ), .C(
        \register[30][25] ), .D(\register[31][25] ), .S0(n1910), .S1(n1869), 
        .Y(n1757) );
  MXI2X1 U1951 ( .A(n1545), .B(n1546), .S0(n1815), .Y(ReadData2_o[26]) );
  MX4X1 U1952 ( .A(n1768), .B(n1766), .C(n1767), .D(n1765), .S0(n1823), .S1(
        n1831), .Y(n1546) );
  MX4X1 U1953 ( .A(n1772), .B(n1770), .C(n1771), .D(n1769), .S0(n1823), .S1(
        n1831), .Y(n1545) );
  MXI4X1 U1954 ( .A(\register[28][26] ), .B(\register[29][26] ), .C(
        \register[30][26] ), .D(\register[31][26] ), .S0(n1911), .S1(n1870), 
        .Y(n1765) );
  MXI2X1 U1955 ( .A(n1547), .B(n1548), .S0(n1815), .Y(ReadData2_o[27]) );
  MX4X1 U1956 ( .A(n1776), .B(n1774), .C(n1775), .D(n1773), .S0(n1823), .S1(
        n1831), .Y(n1548) );
  MX4X1 U1957 ( .A(n1780), .B(n1778), .C(n1779), .D(n1777), .S0(n1823), .S1(
        n1831), .Y(n1547) );
  MXI4X1 U1958 ( .A(\register[28][27] ), .B(\register[29][27] ), .C(
        \register[30][27] ), .D(\register[31][27] ), .S0(n1911), .S1(n1870), 
        .Y(n1773) );
  MXI2X1 U1959 ( .A(n1549), .B(n1550), .S0(n1815), .Y(ReadData2_o[28]) );
  MX4X1 U1960 ( .A(n1784), .B(n1782), .C(n1783), .D(n1781), .S0(n1823), .S1(
        n1831), .Y(n1550) );
  MX4X1 U1961 ( .A(n1788), .B(n1786), .C(n1787), .D(n1785), .S0(n1823), .S1(
        n1831), .Y(n1549) );
  MXI4X1 U1962 ( .A(\register[28][28] ), .B(\register[29][28] ), .C(
        \register[30][28] ), .D(\register[31][28] ), .S0(n1912), .S1(n1871), 
        .Y(n1781) );
  MXI2X1 U1963 ( .A(n1551), .B(n1552), .S0(n1815), .Y(ReadData2_o[29]) );
  MX4X1 U1964 ( .A(n1792), .B(n1790), .C(n1791), .D(n1789), .S0(n1823), .S1(
        n1831), .Y(n1552) );
  MX4X1 U1965 ( .A(n1796), .B(n1794), .C(n1795), .D(n1793), .S0(n1823), .S1(
        n1831), .Y(n1551) );
  MXI4X1 U1966 ( .A(\register[28][29] ), .B(\register[29][29] ), .C(
        \register[30][29] ), .D(\register[31][29] ), .S0(n1913), .S1(n1872), 
        .Y(n1789) );
  MXI2X1 U1967 ( .A(n1553), .B(n1554), .S0(n1815), .Y(ReadData2_o[30]) );
  MX4X1 U1968 ( .A(n1800), .B(n1798), .C(n1799), .D(n1797), .S0(n1823), .S1(
        n1831), .Y(n1554) );
  MX4X1 U1969 ( .A(n1804), .B(n1802), .C(n1803), .D(n1801), .S0(n1823), .S1(
        n1831), .Y(n1553) );
  MXI4X1 U1970 ( .A(\register[28][30] ), .B(\register[29][30] ), .C(
        \register[30][30] ), .D(\register[31][30] ), .S0(n1913), .S1(n1872), 
        .Y(n1797) );
  MXI2X1 U1971 ( .A(n1555), .B(n1556), .S0(n1815), .Y(ReadData2_o[31]) );
  MX4X1 U1972 ( .A(n1808), .B(n1806), .C(n1807), .D(n1805), .S0(n1823), .S1(
        n1831), .Y(n1556) );
  MX4X1 U1973 ( .A(n1812), .B(n1810), .C(n1811), .D(n1809), .S0(n1823), .S1(
        n1831), .Y(n1555) );
  MXI4X1 U1974 ( .A(\register[28][31] ), .B(\register[29][31] ), .C(
        \register[30][31] ), .D(\register[31][31] ), .S0(n1914), .S1(n1873), 
        .Y(n1805) );
  MXI4X1 U1975 ( .A(\register[4][9] ), .B(\register[5][9] ), .C(
        \register[6][9] ), .D(\register[7][9] ), .S0(n1900), .S1(n1859), .Y(
        n1635) );
  MXI4X1 U1976 ( .A(\register[20][9] ), .B(\register[21][9] ), .C(
        \register[22][9] ), .D(\register[23][9] ), .S0(n1899), .S1(n1858), .Y(
        n1631) );
  MXI4X1 U1977 ( .A(\register[4][10] ), .B(\register[5][10] ), .C(
        \register[6][10] ), .D(\register[7][10] ), .S0(n1900), .S1(n1859), .Y(
        n1643) );
  MXI4X1 U1978 ( .A(\register[20][10] ), .B(\register[21][10] ), .C(
        \register[22][10] ), .D(\register[23][10] ), .S0(n1900), .S1(n1859), 
        .Y(n1639) );
  MXI4X1 U1979 ( .A(\register[4][11] ), .B(\register[5][11] ), .C(
        \register[6][11] ), .D(\register[7][11] ), .S0(n1901), .S1(n1860), .Y(
        n1651) );
  MXI4X1 U1980 ( .A(\register[20][11] ), .B(\register[21][11] ), .C(
        \register[22][11] ), .D(\register[23][11] ), .S0(n1901), .S1(n1860), 
        .Y(n1647) );
  MXI4X1 U1981 ( .A(\register[4][12] ), .B(\register[5][12] ), .C(
        \register[6][12] ), .D(\register[7][12] ), .S0(n1902), .S1(n1861), .Y(
        n1659) );
  MXI4X1 U1982 ( .A(\register[20][12] ), .B(\register[21][12] ), .C(
        \register[22][12] ), .D(\register[23][12] ), .S0(n1901), .S1(n1860), 
        .Y(n1655) );
  MXI4X1 U1983 ( .A(\register[4][13] ), .B(\register[5][13] ), .C(
        \register[6][13] ), .D(\register[7][13] ), .S0(n1902), .S1(n1861), .Y(
        n1667) );
  MXI4X1 U1984 ( .A(\register[20][13] ), .B(\register[21][13] ), .C(
        \register[22][13] ), .D(\register[23][13] ), .S0(n1902), .S1(n1861), 
        .Y(n1663) );
  MXI4X1 U1985 ( .A(\register[4][14] ), .B(\register[5][14] ), .C(
        \register[6][14] ), .D(\register[7][14] ), .S0(n1903), .S1(n1862), .Y(
        n1675) );
  MXI4X1 U1986 ( .A(\register[20][14] ), .B(\register[21][14] ), .C(
        \register[22][14] ), .D(\register[23][14] ), .S0(n1903), .S1(n1862), 
        .Y(n1671) );
  MXI4X1 U1987 ( .A(\register[4][15] ), .B(\register[5][15] ), .C(
        \register[6][15] ), .D(\register[7][15] ), .S0(n1904), .S1(n1863), .Y(
        n1683) );
  MXI4X1 U1988 ( .A(\register[20][15] ), .B(\register[21][15] ), .C(
        \register[22][15] ), .D(\register[23][15] ), .S0(n1903), .S1(n1862), 
        .Y(n1679) );
  MXI4X1 U1989 ( .A(\register[4][16] ), .B(\register[5][16] ), .C(
        \register[6][16] ), .D(\register[7][16] ), .S0(n1904), .S1(n1863), .Y(
        n1691) );
  MXI4X1 U1990 ( .A(\register[20][16] ), .B(\register[21][16] ), .C(
        \register[22][16] ), .D(\register[23][16] ), .S0(n1904), .S1(n1863), 
        .Y(n1687) );
  MXI4X1 U1991 ( .A(\register[4][17] ), .B(\register[5][17] ), .C(
        \register[6][17] ), .D(\register[7][17] ), .S0(n1905), .S1(n1864), .Y(
        n1699) );
  MXI4X1 U1992 ( .A(\register[20][17] ), .B(\register[21][17] ), .C(
        \register[22][17] ), .D(\register[23][17] ), .S0(n1905), .S1(n1864), 
        .Y(n1695) );
  MXI4X1 U1993 ( .A(\register[4][18] ), .B(\register[5][18] ), .C(
        \register[6][18] ), .D(\register[7][18] ), .S0(n1906), .S1(n1865), .Y(
        n1707) );
  MXI4X1 U1994 ( .A(\register[20][18] ), .B(\register[21][18] ), .C(
        \register[22][18] ), .D(\register[23][18] ), .S0(n1905), .S1(n1864), 
        .Y(n1703) );
  MXI4X1 U1995 ( .A(\register[4][19] ), .B(\register[5][19] ), .C(
        \register[6][19] ), .D(\register[7][19] ), .S0(n1906), .S1(n1865), .Y(
        n1715) );
  MXI4X1 U1996 ( .A(\register[20][19] ), .B(\register[21][19] ), .C(
        \register[22][19] ), .D(\register[23][19] ), .S0(n1906), .S1(n1865), 
        .Y(n1711) );
  MXI4X1 U1997 ( .A(\register[4][20] ), .B(\register[5][20] ), .C(
        \register[6][20] ), .D(\register[7][20] ), .S0(n1907), .S1(n1866), .Y(
        n1723) );
  MXI4X1 U1998 ( .A(\register[20][20] ), .B(\register[21][20] ), .C(
        \register[22][20] ), .D(\register[23][20] ), .S0(n1907), .S1(n1866), 
        .Y(n1719) );
  MXI4X1 U1999 ( .A(\register[4][21] ), .B(\register[5][21] ), .C(
        \register[6][21] ), .D(\register[7][21] ), .S0(n1908), .S1(n1867), .Y(
        n1731) );
  MXI4X1 U2000 ( .A(\register[20][21] ), .B(\register[21][21] ), .C(
        \register[22][21] ), .D(\register[23][21] ), .S0(n1907), .S1(n1866), 
        .Y(n1727) );
  MXI4X1 U2001 ( .A(\register[4][22] ), .B(\register[5][22] ), .C(
        \register[6][22] ), .D(\register[7][22] ), .S0(n1908), .S1(n1867), .Y(
        n1739) );
  MXI4X1 U2002 ( .A(\register[20][22] ), .B(\register[21][22] ), .C(
        \register[22][22] ), .D(\register[23][22] ), .S0(n1908), .S1(n1867), 
        .Y(n1735) );
  MXI4X1 U2003 ( .A(\register[4][23] ), .B(\register[5][23] ), .C(
        \register[6][23] ), .D(\register[7][23] ), .S0(n1909), .S1(n1868), .Y(
        n1747) );
  MXI4X1 U2004 ( .A(\register[20][23] ), .B(\register[21][23] ), .C(
        \register[22][23] ), .D(\register[23][23] ), .S0(n1909), .S1(n1868), 
        .Y(n1743) );
  MXI4X1 U2005 ( .A(\register[4][24] ), .B(\register[5][24] ), .C(
        \register[6][24] ), .D(\register[7][24] ), .S0(n1910), .S1(n1869), .Y(
        n1755) );
  MXI4X1 U2006 ( .A(\register[20][24] ), .B(\register[21][24] ), .C(
        \register[22][24] ), .D(\register[23][24] ), .S0(n1909), .S1(n1868), 
        .Y(n1751) );
  MXI4X1 U2007 ( .A(\register[4][25] ), .B(\register[5][25] ), .C(
        \register[6][25] ), .D(\register[7][25] ), .S0(n1910), .S1(n1869), .Y(
        n1763) );
  MXI4X1 U2008 ( .A(\register[20][25] ), .B(\register[21][25] ), .C(
        \register[22][25] ), .D(\register[23][25] ), .S0(n1910), .S1(n1869), 
        .Y(n1759) );
  MXI4X1 U2009 ( .A(\register[4][26] ), .B(\register[5][26] ), .C(
        \register[6][26] ), .D(\register[7][26] ), .S0(n1911), .S1(n1870), .Y(
        n1771) );
  MXI4X1 U2010 ( .A(\register[20][26] ), .B(\register[21][26] ), .C(
        \register[22][26] ), .D(\register[23][26] ), .S0(n1911), .S1(n1870), 
        .Y(n1767) );
  MXI4X1 U2011 ( .A(\register[4][27] ), .B(\register[5][27] ), .C(
        \register[6][27] ), .D(\register[7][27] ), .S0(n1912), .S1(n1871), .Y(
        n1779) );
  MXI4X1 U2012 ( .A(\register[20][27] ), .B(\register[21][27] ), .C(
        \register[22][27] ), .D(\register[23][27] ), .S0(n1911), .S1(n1870), 
        .Y(n1775) );
  MXI4X1 U2013 ( .A(\register[4][28] ), .B(\register[5][28] ), .C(
        \register[6][28] ), .D(\register[7][28] ), .S0(n1912), .S1(n1871), .Y(
        n1787) );
  MXI4X1 U2014 ( .A(\register[20][28] ), .B(\register[21][28] ), .C(
        \register[22][28] ), .D(\register[23][28] ), .S0(n1912), .S1(n1871), 
        .Y(n1783) );
  MXI4X1 U2015 ( .A(\register[4][29] ), .B(\register[5][29] ), .C(
        \register[6][29] ), .D(\register[7][29] ), .S0(n1913), .S1(n1872), .Y(
        n1795) );
  MXI4X1 U2016 ( .A(\register[20][29] ), .B(\register[21][29] ), .C(
        \register[22][29] ), .D(\register[23][29] ), .S0(n1913), .S1(n1872), 
        .Y(n1791) );
  MXI4X1 U2017 ( .A(\register[4][30] ), .B(\register[5][30] ), .C(
        \register[6][30] ), .D(\register[7][30] ), .S0(n1914), .S1(n1873), .Y(
        n1803) );
  MXI4X1 U2018 ( .A(\register[20][30] ), .B(\register[21][30] ), .C(
        \register[22][30] ), .D(\register[23][30] ), .S0(n1913), .S1(n1872), 
        .Y(n1799) );
  MXI4X1 U2019 ( .A(\register[4][31] ), .B(\register[5][31] ), .C(
        \register[6][31] ), .D(\register[7][31] ), .S0(n1914), .S1(n1873), .Y(
        n1811) );
  MXI4X1 U2020 ( .A(\register[20][31] ), .B(\register[21][31] ), .C(
        \register[22][31] ), .D(\register[23][31] ), .S0(n1914), .S1(n1873), 
        .Y(n1807) );
  MXI4X1 U2021 ( .A(\register[0][9] ), .B(\register[1][9] ), .C(
        \register[2][9] ), .D(\register[3][9] ), .S0(n1900), .S1(n1859), .Y(
        n1636) );
  MXI4X1 U2022 ( .A(\register[16][9] ), .B(\register[17][9] ), .C(
        \register[18][9] ), .D(\register[19][9] ), .S0(n1899), .S1(n1858), .Y(
        n1632) );
  MXI4X1 U2023 ( .A(\register[0][10] ), .B(\register[1][10] ), .C(
        \register[2][10] ), .D(\register[3][10] ), .S0(n1900), .S1(n1859), .Y(
        n1644) );
  MXI4X1 U2024 ( .A(\register[16][10] ), .B(\register[17][10] ), .C(
        \register[18][10] ), .D(\register[19][10] ), .S0(n1900), .S1(n1859), 
        .Y(n1640) );
  MXI4X1 U2025 ( .A(\register[0][11] ), .B(\register[1][11] ), .C(
        \register[2][11] ), .D(\register[3][11] ), .S0(n1901), .S1(n1860), .Y(
        n1652) );
  MXI4X1 U2026 ( .A(\register[16][11] ), .B(\register[17][11] ), .C(
        \register[18][11] ), .D(\register[19][11] ), .S0(n1901), .S1(n1860), 
        .Y(n1648) );
  MXI4X1 U2027 ( .A(\register[0][12] ), .B(\register[1][12] ), .C(
        \register[2][12] ), .D(\register[3][12] ), .S0(n1902), .S1(n1861), .Y(
        n1660) );
  MXI4X1 U2028 ( .A(\register[16][12] ), .B(\register[17][12] ), .C(
        \register[18][12] ), .D(\register[19][12] ), .S0(n1901), .S1(n1860), 
        .Y(n1656) );
  MXI4X1 U2029 ( .A(\register[0][13] ), .B(\register[1][13] ), .C(
        \register[2][13] ), .D(\register[3][13] ), .S0(n1902), .S1(n1861), .Y(
        n1668) );
  MXI4X1 U2030 ( .A(\register[16][13] ), .B(\register[17][13] ), .C(
        \register[18][13] ), .D(\register[19][13] ), .S0(n1902), .S1(n1861), 
        .Y(n1664) );
  MXI4X1 U2031 ( .A(\register[0][14] ), .B(\register[1][14] ), .C(
        \register[2][14] ), .D(\register[3][14] ), .S0(n1903), .S1(n1862), .Y(
        n1676) );
  MXI4X1 U2032 ( .A(\register[16][14] ), .B(\register[17][14] ), .C(
        \register[18][14] ), .D(\register[19][14] ), .S0(n1903), .S1(n1862), 
        .Y(n1672) );
  MXI4X1 U2033 ( .A(\register[0][15] ), .B(\register[1][15] ), .C(
        \register[2][15] ), .D(\register[3][15] ), .S0(n1904), .S1(n1863), .Y(
        n1684) );
  MXI4X1 U2034 ( .A(\register[16][15] ), .B(\register[17][15] ), .C(
        \register[18][15] ), .D(\register[19][15] ), .S0(n1903), .S1(n1862), 
        .Y(n1680) );
  MXI4X1 U2035 ( .A(\register[0][16] ), .B(\register[1][16] ), .C(
        \register[2][16] ), .D(\register[3][16] ), .S0(n1904), .S1(n1863), .Y(
        n1692) );
  MXI4X1 U2036 ( .A(\register[16][16] ), .B(\register[17][16] ), .C(
        \register[18][16] ), .D(\register[19][16] ), .S0(n1904), .S1(n1863), 
        .Y(n1688) );
  MXI4X1 U2037 ( .A(\register[0][17] ), .B(\register[1][17] ), .C(
        \register[2][17] ), .D(\register[3][17] ), .S0(n1905), .S1(n1864), .Y(
        n1700) );
  MXI4X1 U2038 ( .A(\register[16][17] ), .B(\register[17][17] ), .C(
        \register[18][17] ), .D(\register[19][17] ), .S0(n1905), .S1(n1864), 
        .Y(n1696) );
  MXI4X1 U2039 ( .A(\register[0][18] ), .B(\register[1][18] ), .C(
        \register[2][18] ), .D(\register[3][18] ), .S0(n1906), .S1(n1865), .Y(
        n1708) );
  MXI4X1 U2040 ( .A(\register[16][18] ), .B(\register[17][18] ), .C(
        \register[18][18] ), .D(\register[19][18] ), .S0(n1905), .S1(n1864), 
        .Y(n1704) );
  MXI4X1 U2041 ( .A(\register[0][19] ), .B(\register[1][19] ), .C(
        \register[2][19] ), .D(\register[3][19] ), .S0(n1906), .S1(n1865), .Y(
        n1716) );
  MXI4X1 U2042 ( .A(\register[16][19] ), .B(\register[17][19] ), .C(
        \register[18][19] ), .D(\register[19][19] ), .S0(n1906), .S1(n1865), 
        .Y(n1712) );
  MXI4X1 U2043 ( .A(\register[0][20] ), .B(\register[1][20] ), .C(
        \register[2][20] ), .D(\register[3][20] ), .S0(n1907), .S1(n1866), .Y(
        n1724) );
  MXI4X1 U2044 ( .A(\register[16][20] ), .B(\register[17][20] ), .C(
        \register[18][20] ), .D(\register[19][20] ), .S0(n1907), .S1(n1866), 
        .Y(n1720) );
  MXI4X1 U2045 ( .A(\register[0][21] ), .B(\register[1][21] ), .C(
        \register[2][21] ), .D(\register[3][21] ), .S0(n1908), .S1(n1867), .Y(
        n1732) );
  MXI4X1 U2046 ( .A(\register[16][21] ), .B(\register[17][21] ), .C(
        \register[18][21] ), .D(\register[19][21] ), .S0(n1907), .S1(n1866), 
        .Y(n1728) );
  MXI4X1 U2047 ( .A(\register[0][22] ), .B(\register[1][22] ), .C(
        \register[2][22] ), .D(\register[3][22] ), .S0(n1908), .S1(n1867), .Y(
        n1740) );
  MXI4X1 U2048 ( .A(\register[16][22] ), .B(\register[17][22] ), .C(
        \register[18][22] ), .D(\register[19][22] ), .S0(n1908), .S1(n1867), 
        .Y(n1736) );
  MXI4X1 U2049 ( .A(\register[0][23] ), .B(\register[1][23] ), .C(
        \register[2][23] ), .D(\register[3][23] ), .S0(n1909), .S1(n1868), .Y(
        n1748) );
  MXI4X1 U2050 ( .A(\register[16][23] ), .B(\register[17][23] ), .C(
        \register[18][23] ), .D(\register[19][23] ), .S0(n1909), .S1(n1868), 
        .Y(n1744) );
  MXI4X1 U2051 ( .A(\register[0][24] ), .B(\register[1][24] ), .C(
        \register[2][24] ), .D(\register[3][24] ), .S0(n1910), .S1(n1869), .Y(
        n1756) );
  MXI4X1 U2052 ( .A(\register[16][24] ), .B(\register[17][24] ), .C(
        \register[18][24] ), .D(\register[19][24] ), .S0(n1909), .S1(n1868), 
        .Y(n1752) );
  MXI4X1 U2053 ( .A(\register[0][25] ), .B(\register[1][25] ), .C(
        \register[2][25] ), .D(\register[3][25] ), .S0(n1910), .S1(n1869), .Y(
        n1764) );
  MXI4X1 U2054 ( .A(\register[16][25] ), .B(\register[17][25] ), .C(
        \register[18][25] ), .D(\register[19][25] ), .S0(n1910), .S1(n1869), 
        .Y(n1760) );
  MXI4X1 U2055 ( .A(\register[0][26] ), .B(\register[1][26] ), .C(
        \register[2][26] ), .D(\register[3][26] ), .S0(n1911), .S1(n1870), .Y(
        n1772) );
  MXI4X1 U2056 ( .A(\register[16][26] ), .B(\register[17][26] ), .C(
        \register[18][26] ), .D(\register[19][26] ), .S0(n1911), .S1(n1870), 
        .Y(n1768) );
  MXI4X1 U2057 ( .A(\register[0][27] ), .B(\register[1][27] ), .C(
        \register[2][27] ), .D(\register[3][27] ), .S0(n1912), .S1(n1871), .Y(
        n1780) );
  MXI4X1 U2058 ( .A(\register[16][27] ), .B(\register[17][27] ), .C(
        \register[18][27] ), .D(\register[19][27] ), .S0(n1911), .S1(n1870), 
        .Y(n1776) );
  MXI4X1 U2059 ( .A(\register[0][28] ), .B(\register[1][28] ), .C(
        \register[2][28] ), .D(\register[3][28] ), .S0(n1912), .S1(n1871), .Y(
        n1788) );
  MXI4X1 U2060 ( .A(\register[16][28] ), .B(\register[17][28] ), .C(
        \register[18][28] ), .D(\register[19][28] ), .S0(n1912), .S1(n1871), 
        .Y(n1784) );
  MXI4X1 U2061 ( .A(\register[0][29] ), .B(\register[1][29] ), .C(
        \register[2][29] ), .D(\register[3][29] ), .S0(n1913), .S1(n1872), .Y(
        n1796) );
  MXI4X1 U2062 ( .A(\register[16][29] ), .B(\register[17][29] ), .C(
        \register[18][29] ), .D(\register[19][29] ), .S0(n1913), .S1(n1872), 
        .Y(n1792) );
  MXI4X1 U2063 ( .A(\register[0][30] ), .B(\register[1][30] ), .C(
        \register[2][30] ), .D(\register[3][30] ), .S0(n1914), .S1(n1873), .Y(
        n1804) );
  MXI4X1 U2064 ( .A(\register[16][30] ), .B(\register[17][30] ), .C(
        \register[18][30] ), .D(\register[19][30] ), .S0(n1913), .S1(n1872), 
        .Y(n1800) );
  MXI4X1 U2065 ( .A(\register[0][31] ), .B(\register[1][31] ), .C(
        \register[2][31] ), .D(\register[3][31] ), .S0(n1914), .S1(n1873), .Y(
        n1812) );
  MXI4X1 U2066 ( .A(\register[16][31] ), .B(\register[17][31] ), .C(
        \register[18][31] ), .D(\register[19][31] ), .S0(n1914), .S1(n1873), 
        .Y(n1808) );
  MXI4X1 U2067 ( .A(\register[12][9] ), .B(\register[13][9] ), .C(
        \register[14][9] ), .D(\register[15][9] ), .S0(n1900), .S1(n1859), .Y(
        n1633) );
  MXI4X1 U2068 ( .A(\register[12][10] ), .B(\register[13][10] ), .C(
        \register[14][10] ), .D(\register[15][10] ), .S0(n1900), .S1(n1859), 
        .Y(n1641) );
  MXI4X1 U2069 ( .A(\register[12][11] ), .B(\register[13][11] ), .C(
        \register[14][11] ), .D(\register[15][11] ), .S0(n1901), .S1(n1860), 
        .Y(n1649) );
  MXI4X1 U2070 ( .A(\register[12][12] ), .B(\register[13][12] ), .C(
        \register[14][12] ), .D(\register[15][12] ), .S0(n1902), .S1(n1861), 
        .Y(n1657) );
  MXI4X1 U2071 ( .A(\register[12][13] ), .B(\register[13][13] ), .C(
        \register[14][13] ), .D(\register[15][13] ), .S0(n1902), .S1(n1861), 
        .Y(n1665) );
  MXI4X1 U2072 ( .A(\register[12][14] ), .B(\register[13][14] ), .C(
        \register[14][14] ), .D(\register[15][14] ), .S0(n1903), .S1(n1862), 
        .Y(n1673) );
  MXI4X1 U2073 ( .A(\register[12][15] ), .B(\register[13][15] ), .C(
        \register[14][15] ), .D(\register[15][15] ), .S0(n1904), .S1(n1863), 
        .Y(n1681) );
  MXI4X1 U2074 ( .A(\register[12][16] ), .B(\register[13][16] ), .C(
        \register[14][16] ), .D(\register[15][16] ), .S0(n1904), .S1(n1863), 
        .Y(n1689) );
  MXI4X1 U2075 ( .A(\register[12][17] ), .B(\register[13][17] ), .C(
        \register[14][17] ), .D(\register[15][17] ), .S0(n1905), .S1(n1864), 
        .Y(n1697) );
  MXI4X1 U2076 ( .A(\register[12][18] ), .B(\register[13][18] ), .C(
        \register[14][18] ), .D(\register[15][18] ), .S0(n1906), .S1(n1865), 
        .Y(n1705) );
  MXI4X1 U2077 ( .A(\register[12][19] ), .B(\register[13][19] ), .C(
        \register[14][19] ), .D(\register[15][19] ), .S0(n1906), .S1(n1865), 
        .Y(n1713) );
  MXI4X1 U2078 ( .A(\register[12][20] ), .B(\register[13][20] ), .C(
        \register[14][20] ), .D(\register[15][20] ), .S0(n1907), .S1(n1866), 
        .Y(n1721) );
  MXI4X1 U2079 ( .A(\register[12][21] ), .B(\register[13][21] ), .C(
        \register[14][21] ), .D(\register[15][21] ), .S0(n1908), .S1(n1867), 
        .Y(n1729) );
  MXI4X1 U2080 ( .A(\register[12][22] ), .B(\register[13][22] ), .C(
        \register[14][22] ), .D(\register[15][22] ), .S0(n1908), .S1(n1867), 
        .Y(n1737) );
  MXI4X1 U2081 ( .A(\register[12][23] ), .B(\register[13][23] ), .C(
        \register[14][23] ), .D(\register[15][23] ), .S0(n1909), .S1(n1868), 
        .Y(n1745) );
  MXI4X1 U2082 ( .A(\register[12][24] ), .B(\register[13][24] ), .C(
        \register[14][24] ), .D(\register[15][24] ), .S0(n1910), .S1(n1869), 
        .Y(n1753) );
  MXI4X1 U2083 ( .A(\register[12][25] ), .B(\register[13][25] ), .C(
        \register[14][25] ), .D(\register[15][25] ), .S0(n1910), .S1(n1869), 
        .Y(n1761) );
  MXI4X1 U2084 ( .A(\register[12][26] ), .B(\register[13][26] ), .C(
        \register[14][26] ), .D(\register[15][26] ), .S0(n1911), .S1(n1870), 
        .Y(n1769) );
  MXI4X1 U2085 ( .A(\register[12][27] ), .B(\register[13][27] ), .C(
        \register[14][27] ), .D(\register[15][27] ), .S0(n1912), .S1(n1871), 
        .Y(n1777) );
  MXI4X1 U2086 ( .A(\register[12][28] ), .B(\register[13][28] ), .C(
        \register[14][28] ), .D(\register[15][28] ), .S0(n1912), .S1(n1871), 
        .Y(n1785) );
  MXI4X1 U2087 ( .A(\register[12][29] ), .B(\register[13][29] ), .C(
        \register[14][29] ), .D(\register[15][29] ), .S0(n1913), .S1(n1872), 
        .Y(n1793) );
  MXI4X1 U2088 ( .A(\register[12][30] ), .B(\register[13][30] ), .C(
        \register[14][30] ), .D(\register[15][30] ), .S0(n1914), .S1(n1873), 
        .Y(n1801) );
  MXI4X1 U2089 ( .A(\register[12][31] ), .B(\register[13][31] ), .C(
        \register[14][31] ), .D(\register[15][31] ), .S0(n1914), .S1(n1873), 
        .Y(n1809) );
  MXI4X1 U2090 ( .A(\register[8][9] ), .B(\register[9][9] ), .C(
        \register[10][9] ), .D(\register[11][9] ), .S0(n1900), .S1(n1859), .Y(
        n1634) );
  MXI4X1 U2091 ( .A(\register[24][9] ), .B(\register[25][9] ), .C(
        \register[26][9] ), .D(\register[27][9] ), .S0(n1899), .S1(n1858), .Y(
        n1630) );
  MXI4X1 U2092 ( .A(\register[8][10] ), .B(\register[9][10] ), .C(
        \register[10][10] ), .D(\register[11][10] ), .S0(n1900), .S1(n1859), 
        .Y(n1642) );
  MXI4X1 U2093 ( .A(\register[24][10] ), .B(\register[25][10] ), .C(
        \register[26][10] ), .D(\register[27][10] ), .S0(n1900), .S1(n1859), 
        .Y(n1638) );
  MXI4X1 U2094 ( .A(\register[8][11] ), .B(\register[9][11] ), .C(
        \register[10][11] ), .D(\register[11][11] ), .S0(n1901), .S1(n1860), 
        .Y(n1650) );
  MXI4X1 U2095 ( .A(\register[24][11] ), .B(\register[25][11] ), .C(
        \register[26][11] ), .D(\register[27][11] ), .S0(n1901), .S1(n1860), 
        .Y(n1646) );
  MXI4X1 U2096 ( .A(\register[8][12] ), .B(\register[9][12] ), .C(
        \register[10][12] ), .D(\register[11][12] ), .S0(n1902), .S1(n1861), 
        .Y(n1658) );
  MXI4X1 U2097 ( .A(\register[24][12] ), .B(\register[25][12] ), .C(
        \register[26][12] ), .D(\register[27][12] ), .S0(n1901), .S1(n1860), 
        .Y(n1654) );
  MXI4X1 U2098 ( .A(\register[8][13] ), .B(\register[9][13] ), .C(
        \register[10][13] ), .D(\register[11][13] ), .S0(n1902), .S1(n1861), 
        .Y(n1666) );
  MXI4X1 U2099 ( .A(\register[24][13] ), .B(\register[25][13] ), .C(
        \register[26][13] ), .D(\register[27][13] ), .S0(n1902), .S1(n1861), 
        .Y(n1662) );
  MXI4X1 U2100 ( .A(\register[8][14] ), .B(\register[9][14] ), .C(
        \register[10][14] ), .D(\register[11][14] ), .S0(n1903), .S1(n1862), 
        .Y(n1674) );
  MXI4X1 U2101 ( .A(\register[24][14] ), .B(\register[25][14] ), .C(
        \register[26][14] ), .D(\register[27][14] ), .S0(n1903), .S1(n1862), 
        .Y(n1670) );
  MXI4X1 U2102 ( .A(\register[8][15] ), .B(\register[9][15] ), .C(
        \register[10][15] ), .D(\register[11][15] ), .S0(n1904), .S1(n1863), 
        .Y(n1682) );
  MXI4X1 U2103 ( .A(\register[24][15] ), .B(\register[25][15] ), .C(
        \register[26][15] ), .D(\register[27][15] ), .S0(n1903), .S1(n1862), 
        .Y(n1678) );
  MXI4X1 U2104 ( .A(\register[8][16] ), .B(\register[9][16] ), .C(
        \register[10][16] ), .D(\register[11][16] ), .S0(n1904), .S1(n1863), 
        .Y(n1690) );
  MXI4X1 U2105 ( .A(\register[24][16] ), .B(\register[25][16] ), .C(
        \register[26][16] ), .D(\register[27][16] ), .S0(n1904), .S1(n1863), 
        .Y(n1686) );
  MXI4X1 U2106 ( .A(\register[8][17] ), .B(\register[9][17] ), .C(
        \register[10][17] ), .D(\register[11][17] ), .S0(n1905), .S1(n1864), 
        .Y(n1698) );
  MXI4X1 U2107 ( .A(\register[24][17] ), .B(\register[25][17] ), .C(
        \register[26][17] ), .D(\register[27][17] ), .S0(n1905), .S1(n1864), 
        .Y(n1694) );
  MXI4X1 U2108 ( .A(\register[8][18] ), .B(\register[9][18] ), .C(
        \register[10][18] ), .D(\register[11][18] ), .S0(n1906), .S1(n1865), 
        .Y(n1706) );
  MXI4X1 U2109 ( .A(\register[24][18] ), .B(\register[25][18] ), .C(
        \register[26][18] ), .D(\register[27][18] ), .S0(n1905), .S1(n1864), 
        .Y(n1702) );
  MXI4X1 U2110 ( .A(\register[8][19] ), .B(\register[9][19] ), .C(
        \register[10][19] ), .D(\register[11][19] ), .S0(n1906), .S1(n1865), 
        .Y(n1714) );
  MXI4X1 U2111 ( .A(\register[24][19] ), .B(\register[25][19] ), .C(
        \register[26][19] ), .D(\register[27][19] ), .S0(n1906), .S1(n1865), 
        .Y(n1710) );
  MXI4X1 U2112 ( .A(\register[8][20] ), .B(\register[9][20] ), .C(
        \register[10][20] ), .D(\register[11][20] ), .S0(n1907), .S1(n1866), 
        .Y(n1722) );
  MXI4X1 U2113 ( .A(\register[24][20] ), .B(\register[25][20] ), .C(
        \register[26][20] ), .D(\register[27][20] ), .S0(n1907), .S1(n1866), 
        .Y(n1718) );
  MXI4X1 U2114 ( .A(\register[8][21] ), .B(\register[9][21] ), .C(
        \register[10][21] ), .D(\register[11][21] ), .S0(n1908), .S1(n1867), 
        .Y(n1730) );
  MXI4X1 U2115 ( .A(\register[24][21] ), .B(\register[25][21] ), .C(
        \register[26][21] ), .D(\register[27][21] ), .S0(n1907), .S1(n1866), 
        .Y(n1726) );
  MXI4X1 U2116 ( .A(\register[8][22] ), .B(\register[9][22] ), .C(
        \register[10][22] ), .D(\register[11][22] ), .S0(n1908), .S1(n1867), 
        .Y(n1738) );
  MXI4X1 U2117 ( .A(\register[24][22] ), .B(\register[25][22] ), .C(
        \register[26][22] ), .D(\register[27][22] ), .S0(n1908), .S1(n1867), 
        .Y(n1734) );
  MXI4X1 U2118 ( .A(\register[8][23] ), .B(\register[9][23] ), .C(
        \register[10][23] ), .D(\register[11][23] ), .S0(n1909), .S1(n1868), 
        .Y(n1746) );
  MXI4X1 U2119 ( .A(\register[24][23] ), .B(\register[25][23] ), .C(
        \register[26][23] ), .D(\register[27][23] ), .S0(n1909), .S1(n1868), 
        .Y(n1742) );
  MXI4X1 U2120 ( .A(\register[8][24] ), .B(\register[9][24] ), .C(
        \register[10][24] ), .D(\register[11][24] ), .S0(n1910), .S1(n1869), 
        .Y(n1754) );
  MXI4X1 U2121 ( .A(\register[24][24] ), .B(\register[25][24] ), .C(
        \register[26][24] ), .D(\register[27][24] ), .S0(n1909), .S1(n1868), 
        .Y(n1750) );
  MXI4X1 U2122 ( .A(\register[8][25] ), .B(\register[9][25] ), .C(
        \register[10][25] ), .D(\register[11][25] ), .S0(n1910), .S1(n1869), 
        .Y(n1762) );
  MXI4X1 U2123 ( .A(\register[24][25] ), .B(\register[25][25] ), .C(
        \register[26][25] ), .D(\register[27][25] ), .S0(n1910), .S1(n1869), 
        .Y(n1758) );
  MXI4X1 U2124 ( .A(\register[8][26] ), .B(\register[9][26] ), .C(
        \register[10][26] ), .D(\register[11][26] ), .S0(n1911), .S1(n1870), 
        .Y(n1770) );
  MXI4X1 U2125 ( .A(\register[24][26] ), .B(\register[25][26] ), .C(
        \register[26][26] ), .D(\register[27][26] ), .S0(n1911), .S1(n1870), 
        .Y(n1766) );
  MXI4X1 U2126 ( .A(\register[8][27] ), .B(\register[9][27] ), .C(
        \register[10][27] ), .D(\register[11][27] ), .S0(n1912), .S1(n1871), 
        .Y(n1778) );
  MXI4X1 U2127 ( .A(\register[24][27] ), .B(\register[25][27] ), .C(
        \register[26][27] ), .D(\register[27][27] ), .S0(n1911), .S1(n1870), 
        .Y(n1774) );
  MXI4X1 U2128 ( .A(\register[8][28] ), .B(\register[9][28] ), .C(
        \register[10][28] ), .D(\register[11][28] ), .S0(n1912), .S1(n1871), 
        .Y(n1786) );
  MXI4X1 U2129 ( .A(\register[24][28] ), .B(\register[25][28] ), .C(
        \register[26][28] ), .D(\register[27][28] ), .S0(n1912), .S1(n1871), 
        .Y(n1782) );
  MXI4X1 U2130 ( .A(\register[8][29] ), .B(\register[9][29] ), .C(
        \register[10][29] ), .D(\register[11][29] ), .S0(n1913), .S1(n1872), 
        .Y(n1794) );
  MXI4X1 U2131 ( .A(\register[24][29] ), .B(\register[25][29] ), .C(
        \register[26][29] ), .D(\register[27][29] ), .S0(n1913), .S1(n1872), 
        .Y(n1790) );
  MXI4X1 U2132 ( .A(\register[8][30] ), .B(\register[9][30] ), .C(
        \register[10][30] ), .D(\register[11][30] ), .S0(n1914), .S1(n1873), 
        .Y(n1802) );
  MXI4X1 U2133 ( .A(\register[24][30] ), .B(\register[25][30] ), .C(
        \register[26][30] ), .D(\register[27][30] ), .S0(n1913), .S1(n1872), 
        .Y(n1798) );
  MXI4X1 U2134 ( .A(\register[8][31] ), .B(\register[9][31] ), .C(
        \register[10][31] ), .D(\register[11][31] ), .S0(n1914), .S1(n1873), 
        .Y(n1810) );
  MXI4X1 U2135 ( .A(\register[24][31] ), .B(\register[25][31] ), .C(
        \register[26][31] ), .D(\register[27][31] ), .S0(n1914), .S1(n1873), 
        .Y(n1806) );
  MX4X1 U2136 ( .A(n1208), .B(n1206), .C(n1207), .D(n1205), .S0(n1396), .S1(
        n1404), .Y(n20) );
  MX4X1 U2137 ( .A(n1212), .B(n1210), .C(n1211), .D(n1209), .S0(n1396), .S1(
        n1404), .Y(n19) );
  MXI4X1 U2138 ( .A(\register[28][9] ), .B(\register[29][9] ), .C(
        \register[30][9] ), .D(\register[31][9] ), .S0(n1475), .S1(n1434), .Y(
        n1205) );
  MX4X1 U2139 ( .A(n1224), .B(n1222), .C(n1223), .D(n1221), .S0(n1396), .S1(
        n1404), .Y(n24) );
  MX4X1 U2140 ( .A(n1228), .B(n1226), .C(n1227), .D(n1225), .S0(n1396), .S1(
        n1404), .Y(n23) );
  MXI4X1 U2141 ( .A(\register[28][11] ), .B(\register[29][11] ), .C(
        \register[30][11] ), .D(\register[31][11] ), .S0(n1477), .S1(n1436), 
        .Y(n1221) );
  MX4X1 U2142 ( .A(n1216), .B(n1214), .C(n1215), .D(n1213), .S0(n1396), .S1(
        n1404), .Y(n22) );
  MX4X1 U2143 ( .A(n1220), .B(n1218), .C(n1219), .D(n1217), .S0(n1396), .S1(
        n1404), .Y(n21) );
  MXI4X1 U2144 ( .A(\register[28][10] ), .B(\register[29][10] ), .C(
        \register[30][10] ), .D(\register[31][10] ), .S0(n1476), .S1(n1435), 
        .Y(n1213) );
  MX4X1 U2145 ( .A(n1232), .B(n1230), .C(n1231), .D(n1229), .S0(n1396), .S1(
        n1404), .Y(n26) );
  MX4X1 U2146 ( .A(n1236), .B(n1234), .C(n1235), .D(n1233), .S0(n1396), .S1(
        n1405), .Y(n25) );
  MXI4X1 U2147 ( .A(\register[28][12] ), .B(\register[29][12] ), .C(
        \register[30][12] ), .D(\register[31][12] ), .S0(n1477), .S1(n1436), 
        .Y(n1229) );
  MXI4X1 U2148 ( .A(\register[4][9] ), .B(\register[5][9] ), .C(
        \register[6][9] ), .D(\register[7][9] ), .S0(n1476), .S1(n1435), .Y(
        n1211) );
  MXI4X1 U2149 ( .A(\register[20][9] ), .B(\register[21][9] ), .C(
        \register[22][9] ), .D(\register[23][9] ), .S0(n1475), .S1(n1434), .Y(
        n1207) );
  MXI4X1 U2150 ( .A(\register[4][10] ), .B(\register[5][10] ), .C(
        \register[6][10] ), .D(\register[7][10] ), .S0(n1476), .S1(n1435), .Y(
        n1219) );
  MXI4X1 U2151 ( .A(\register[20][10] ), .B(\register[21][10] ), .C(
        \register[22][10] ), .D(\register[23][10] ), .S0(n1476), .S1(n1435), 
        .Y(n1215) );
  MXI4X1 U2152 ( .A(\register[4][11] ), .B(\register[5][11] ), .C(
        \register[6][11] ), .D(\register[7][11] ), .S0(n1477), .S1(n1436), .Y(
        n1227) );
  MXI4X1 U2153 ( .A(\register[20][11] ), .B(\register[21][11] ), .C(
        \register[22][11] ), .D(\register[23][11] ), .S0(n1477), .S1(n1436), 
        .Y(n1223) );
  MXI4X1 U2154 ( .A(\register[4][12] ), .B(\register[5][12] ), .C(
        \register[6][12] ), .D(\register[7][12] ), .S0(n1478), .S1(n1437), .Y(
        n1235) );
  MXI4X1 U2155 ( .A(\register[20][12] ), .B(\register[21][12] ), .C(
        \register[22][12] ), .D(\register[23][12] ), .S0(n1477), .S1(n1436), 
        .Y(n1231) );
  MXI4X1 U2156 ( .A(\register[0][9] ), .B(\register[1][9] ), .C(
        \register[2][9] ), .D(\register[3][9] ), .S0(n1476), .S1(n1435), .Y(
        n1212) );
  MXI4X1 U2157 ( .A(\register[16][9] ), .B(\register[17][9] ), .C(
        \register[18][9] ), .D(\register[19][9] ), .S0(n1475), .S1(n1434), .Y(
        n1208) );
  MXI4X1 U2158 ( .A(\register[0][10] ), .B(\register[1][10] ), .C(
        \register[2][10] ), .D(\register[3][10] ), .S0(n1476), .S1(n1435), .Y(
        n1220) );
  MXI4X1 U2159 ( .A(\register[16][10] ), .B(\register[17][10] ), .C(
        \register[18][10] ), .D(\register[19][10] ), .S0(n1476), .S1(n1435), 
        .Y(n1216) );
  MXI4X1 U2160 ( .A(\register[0][11] ), .B(\register[1][11] ), .C(
        \register[2][11] ), .D(\register[3][11] ), .S0(n1477), .S1(n1436), .Y(
        n1228) );
  MXI4X1 U2161 ( .A(\register[16][11] ), .B(\register[17][11] ), .C(
        \register[18][11] ), .D(\register[19][11] ), .S0(n1477), .S1(n1436), 
        .Y(n1224) );
  MXI4X1 U2162 ( .A(\register[0][12] ), .B(\register[1][12] ), .C(
        \register[2][12] ), .D(\register[3][12] ), .S0(n1478), .S1(n1437), .Y(
        n1236) );
  MXI4X1 U2163 ( .A(\register[16][12] ), .B(\register[17][12] ), .C(
        \register[18][12] ), .D(\register[19][12] ), .S0(n1477), .S1(n1436), 
        .Y(n1232) );
  MXI4X1 U2164 ( .A(\register[12][9] ), .B(\register[13][9] ), .C(
        \register[14][9] ), .D(\register[15][9] ), .S0(n1476), .S1(n1435), .Y(
        n1209) );
  MXI4X1 U2165 ( .A(\register[12][10] ), .B(\register[13][10] ), .C(
        \register[14][10] ), .D(\register[15][10] ), .S0(n1476), .S1(n1435), 
        .Y(n1217) );
  MXI4X1 U2166 ( .A(\register[12][11] ), .B(\register[13][11] ), .C(
        \register[14][11] ), .D(\register[15][11] ), .S0(n1477), .S1(n1436), 
        .Y(n1225) );
  MXI4X1 U2167 ( .A(\register[12][12] ), .B(\register[13][12] ), .C(
        \register[14][12] ), .D(\register[15][12] ), .S0(n1478), .S1(n1437), 
        .Y(n1233) );
  MXI4X1 U2168 ( .A(\register[8][9] ), .B(\register[9][9] ), .C(
        \register[10][9] ), .D(\register[11][9] ), .S0(n1476), .S1(n1435), .Y(
        n1210) );
  MXI4X1 U2169 ( .A(\register[24][9] ), .B(\register[25][9] ), .C(
        \register[26][9] ), .D(\register[27][9] ), .S0(n1475), .S1(n1434), .Y(
        n1206) );
  MXI4X1 U2170 ( .A(\register[8][10] ), .B(\register[9][10] ), .C(
        \register[10][10] ), .D(\register[11][10] ), .S0(n1476), .S1(n1435), 
        .Y(n1218) );
  MXI4X1 U2171 ( .A(\register[24][10] ), .B(\register[25][10] ), .C(
        \register[26][10] ), .D(\register[27][10] ), .S0(n1476), .S1(n1435), 
        .Y(n1214) );
  MXI4X1 U2172 ( .A(\register[8][11] ), .B(\register[9][11] ), .C(
        \register[10][11] ), .D(\register[11][11] ), .S0(n1477), .S1(n1436), 
        .Y(n1226) );
  MXI4X1 U2173 ( .A(\register[24][11] ), .B(\register[25][11] ), .C(
        \register[26][11] ), .D(\register[27][11] ), .S0(n1477), .S1(n1436), 
        .Y(n1222) );
  MXI4X1 U2174 ( .A(\register[8][12] ), .B(\register[9][12] ), .C(
        \register[10][12] ), .D(\register[11][12] ), .S0(n1478), .S1(n1437), 
        .Y(n1234) );
  MXI4X1 U2175 ( .A(\register[24][12] ), .B(\register[25][12] ), .C(
        \register[26][12] ), .D(\register[27][12] ), .S0(n1477), .S1(n1436), 
        .Y(n1230) );
  MX4X1 U2176 ( .A(n1248), .B(n1246), .C(n1247), .D(n1245), .S0(n1397), .S1(
        n1405), .Y(n30) );
  MX4X1 U2177 ( .A(n1252), .B(n1250), .C(n1251), .D(n1249), .S0(n1397), .S1(
        n1405), .Y(n29) );
  MXI4X1 U2178 ( .A(\register[28][14] ), .B(\register[29][14] ), .C(
        \register[30][14] ), .D(\register[31][14] ), .S0(n1479), .S1(n1438), 
        .Y(n1245) );
  MX4X1 U2179 ( .A(n1264), .B(n1262), .C(n1263), .D(n1261), .S0(n1397), .S1(
        n1405), .Y(n34) );
  MX4X1 U2180 ( .A(n1268), .B(n1266), .C(n1267), .D(n1265), .S0(n1397), .S1(
        n1405), .Y(n33) );
  MXI4X1 U2181 ( .A(\register[28][16] ), .B(\register[29][16] ), .C(
        \register[30][16] ), .D(\register[31][16] ), .S0(n1480), .S1(n1439), 
        .Y(n1261) );
  MX4X1 U2182 ( .A(n1272), .B(n1270), .C(n1271), .D(n1269), .S0(n1397), .S1(
        n1405), .Y(n36) );
  MX4X1 U2183 ( .A(n1276), .B(n1274), .C(n1275), .D(n1273), .S0(n1397), .S1(
        n1405), .Y(n35) );
  MXI4X1 U2184 ( .A(\register[28][17] ), .B(\register[29][17] ), .C(
        \register[30][17] ), .D(\register[31][17] ), .S0(n1481), .S1(n1440), 
        .Y(n1269) );
  MX4X1 U2185 ( .A(n1288), .B(n1286), .C(n1287), .D(n1285), .S0(n1397), .S1(
        n1406), .Y(n1108) );
  MX4X1 U2186 ( .A(n1292), .B(n1290), .C(n1291), .D(n1289), .S0(n1397), .S1(
        n1406), .Y(n1107) );
  MXI4X1 U2187 ( .A(\register[28][19] ), .B(\register[29][19] ), .C(
        \register[30][19] ), .D(\register[31][19] ), .S0(n1482), .S1(n1441), 
        .Y(n1285) );
  MX4X1 U2188 ( .A(n1240), .B(n1238), .C(n1239), .D(n1237), .S0(n1396), .S1(
        n1405), .Y(n28) );
  MX4X1 U2189 ( .A(n1244), .B(n1242), .C(n1243), .D(n1241), .S0(n1396), .S1(
        n1405), .Y(n27) );
  MXI4X1 U2190 ( .A(\register[28][13] ), .B(\register[29][13] ), .C(
        \register[30][13] ), .D(\register[31][13] ), .S0(n1478), .S1(n1437), 
        .Y(n1237) );
  MX4X1 U2191 ( .A(n1304), .B(n1302), .C(n1303), .D(n1301), .S0(n1398), .S1(
        n1406), .Y(n1112) );
  MX4X1 U2192 ( .A(n1308), .B(n1306), .C(n1307), .D(n1305), .S0(n1398), .S1(
        n1406), .Y(n1111) );
  MXI4X1 U2193 ( .A(\register[28][21] ), .B(\register[29][21] ), .C(
        \register[30][21] ), .D(\register[31][21] ), .S0(n1483), .S1(n1442), 
        .Y(n1301) );
  MX4X1 U2194 ( .A(n1296), .B(n1294), .C(n1295), .D(n1293), .S0(n1398), .S1(
        n1406), .Y(n1110) );
  MX4X1 U2195 ( .A(n1300), .B(n1298), .C(n1299), .D(n1297), .S0(n1398), .S1(
        n1406), .Y(n1109) );
  MXI4X1 U2196 ( .A(\register[28][20] ), .B(\register[29][20] ), .C(
        \register[30][20] ), .D(\register[31][20] ), .S0(n1483), .S1(n1442), 
        .Y(n1293) );
  MX4X1 U2197 ( .A(n1280), .B(n1278), .C(n1279), .D(n1277), .S0(n1397), .S1(
        n1405), .Y(n1106) );
  MX4X1 U2198 ( .A(n1284), .B(n1282), .C(n1283), .D(n1281), .S0(n1397), .S1(
        n1405), .Y(n37) );
  MXI4X1 U2199 ( .A(\register[28][18] ), .B(\register[29][18] ), .C(
        \register[30][18] ), .D(\register[31][18] ), .S0(n1481), .S1(n1440), 
        .Y(n1277) );
  MX4X1 U2200 ( .A(n1256), .B(n1254), .C(n1255), .D(n1253), .S0(n1397), .S1(
        n1405), .Y(n32) );
  MX4X1 U2201 ( .A(n1260), .B(n1258), .C(n1259), .D(n1257), .S0(n1397), .S1(
        n1405), .Y(n31) );
  MXI4X1 U2202 ( .A(\register[28][15] ), .B(\register[29][15] ), .C(
        \register[30][15] ), .D(\register[31][15] ), .S0(n1479), .S1(n1438), 
        .Y(n1253) );
  MXI4X1 U2203 ( .A(\register[4][13] ), .B(\register[5][13] ), .C(
        \register[6][13] ), .D(\register[7][13] ), .S0(n1478), .S1(n1437), .Y(
        n1243) );
  MXI4X1 U2204 ( .A(\register[20][13] ), .B(\register[21][13] ), .C(
        \register[22][13] ), .D(\register[23][13] ), .S0(n1478), .S1(n1437), 
        .Y(n1239) );
  MXI4X1 U2205 ( .A(\register[4][14] ), .B(\register[5][14] ), .C(
        \register[6][14] ), .D(\register[7][14] ), .S0(n1479), .S1(n1438), .Y(
        n1251) );
  MXI4X1 U2206 ( .A(\register[20][14] ), .B(\register[21][14] ), .C(
        \register[22][14] ), .D(\register[23][14] ), .S0(n1479), .S1(n1438), 
        .Y(n1247) );
  MXI4X1 U2207 ( .A(\register[4][16] ), .B(\register[5][16] ), .C(
        \register[6][16] ), .D(\register[7][16] ), .S0(n1480), .S1(n1439), .Y(
        n1267) );
  MXI4X1 U2208 ( .A(\register[20][16] ), .B(\register[21][16] ), .C(
        \register[22][16] ), .D(\register[23][16] ), .S0(n1480), .S1(n1439), 
        .Y(n1263) );
  MXI4X1 U2209 ( .A(\register[4][15] ), .B(\register[5][15] ), .C(
        \register[6][15] ), .D(\register[7][15] ), .S0(n1480), .S1(n1439), .Y(
        n1259) );
  MXI4X1 U2210 ( .A(\register[20][15] ), .B(\register[21][15] ), .C(
        \register[22][15] ), .D(\register[23][15] ), .S0(n1479), .S1(n1438), 
        .Y(n1255) );
  MXI4X1 U2211 ( .A(\register[4][17] ), .B(\register[5][17] ), .C(
        \register[6][17] ), .D(\register[7][17] ), .S0(n1481), .S1(n1440), .Y(
        n1275) );
  MXI4X1 U2212 ( .A(\register[20][17] ), .B(\register[21][17] ), .C(
        \register[22][17] ), .D(\register[23][17] ), .S0(n1481), .S1(n1440), 
        .Y(n1271) );
  MXI4X1 U2213 ( .A(\register[4][18] ), .B(\register[5][18] ), .C(
        \register[6][18] ), .D(\register[7][18] ), .S0(n1482), .S1(n1441), .Y(
        n1283) );
  MXI4X1 U2214 ( .A(\register[20][18] ), .B(\register[21][18] ), .C(
        \register[22][18] ), .D(\register[23][18] ), .S0(n1481), .S1(n1440), 
        .Y(n1279) );
  MXI4X1 U2215 ( .A(\register[4][19] ), .B(\register[5][19] ), .C(
        \register[6][19] ), .D(\register[7][19] ), .S0(n1482), .S1(n1441), .Y(
        n1291) );
  MXI4X1 U2216 ( .A(\register[20][19] ), .B(\register[21][19] ), .C(
        \register[22][19] ), .D(\register[23][19] ), .S0(n1482), .S1(n1441), 
        .Y(n1287) );
  MXI4X1 U2217 ( .A(\register[4][20] ), .B(\register[5][20] ), .C(
        \register[6][20] ), .D(\register[7][20] ), .S0(n1483), .S1(n1442), .Y(
        n1299) );
  MXI4X1 U2218 ( .A(\register[20][20] ), .B(\register[21][20] ), .C(
        \register[22][20] ), .D(\register[23][20] ), .S0(n1483), .S1(n1442), 
        .Y(n1295) );
  MXI4X1 U2219 ( .A(\register[4][21] ), .B(\register[5][21] ), .C(
        \register[6][21] ), .D(\register[7][21] ), .S0(n1484), .S1(n1443), .Y(
        n1307) );
  MXI4X1 U2220 ( .A(\register[20][21] ), .B(\register[21][21] ), .C(
        \register[22][21] ), .D(\register[23][21] ), .S0(n1483), .S1(n1442), 
        .Y(n1303) );
  MXI4X1 U2221 ( .A(\register[0][13] ), .B(\register[1][13] ), .C(
        \register[2][13] ), .D(\register[3][13] ), .S0(n1478), .S1(n1437), .Y(
        n1244) );
  MXI4X1 U2222 ( .A(\register[16][13] ), .B(\register[17][13] ), .C(
        \register[18][13] ), .D(\register[19][13] ), .S0(n1478), .S1(n1437), 
        .Y(n1240) );
  MXI4X1 U2223 ( .A(\register[0][14] ), .B(\register[1][14] ), .C(
        \register[2][14] ), .D(\register[3][14] ), .S0(n1479), .S1(n1438), .Y(
        n1252) );
  MXI4X1 U2224 ( .A(\register[16][14] ), .B(\register[17][14] ), .C(
        \register[18][14] ), .D(\register[19][14] ), .S0(n1479), .S1(n1438), 
        .Y(n1248) );
  MXI4X1 U2225 ( .A(\register[0][16] ), .B(\register[1][16] ), .C(
        \register[2][16] ), .D(\register[3][16] ), .S0(n1480), .S1(n1439), .Y(
        n1268) );
  MXI4X1 U2226 ( .A(\register[16][16] ), .B(\register[17][16] ), .C(
        \register[18][16] ), .D(\register[19][16] ), .S0(n1480), .S1(n1439), 
        .Y(n1264) );
  MXI4X1 U2227 ( .A(\register[0][15] ), .B(\register[1][15] ), .C(
        \register[2][15] ), .D(\register[3][15] ), .S0(n1480), .S1(n1439), .Y(
        n1260) );
  MXI4X1 U2228 ( .A(\register[16][15] ), .B(\register[17][15] ), .C(
        \register[18][15] ), .D(\register[19][15] ), .S0(n1479), .S1(n1438), 
        .Y(n1256) );
  MXI4X1 U2229 ( .A(\register[0][17] ), .B(\register[1][17] ), .C(
        \register[2][17] ), .D(\register[3][17] ), .S0(n1481), .S1(n1440), .Y(
        n1276) );
  MXI4X1 U2230 ( .A(\register[16][17] ), .B(\register[17][17] ), .C(
        \register[18][17] ), .D(\register[19][17] ), .S0(n1481), .S1(n1440), 
        .Y(n1272) );
  MXI4X1 U2231 ( .A(\register[0][18] ), .B(\register[1][18] ), .C(
        \register[2][18] ), .D(\register[3][18] ), .S0(n1482), .S1(n1441), .Y(
        n1284) );
  MXI4X1 U2232 ( .A(\register[16][18] ), .B(\register[17][18] ), .C(
        \register[18][18] ), .D(\register[19][18] ), .S0(n1481), .S1(n1440), 
        .Y(n1280) );
  MXI4X1 U2233 ( .A(\register[0][19] ), .B(\register[1][19] ), .C(
        \register[2][19] ), .D(\register[3][19] ), .S0(n1482), .S1(n1441), .Y(
        n1292) );
  MXI4X1 U2234 ( .A(\register[16][19] ), .B(\register[17][19] ), .C(
        \register[18][19] ), .D(\register[19][19] ), .S0(n1482), .S1(n1441), 
        .Y(n1288) );
  MXI4X1 U2235 ( .A(\register[0][20] ), .B(\register[1][20] ), .C(
        \register[2][20] ), .D(\register[3][20] ), .S0(n1483), .S1(n1442), .Y(
        n1300) );
  MXI4X1 U2236 ( .A(\register[16][20] ), .B(\register[17][20] ), .C(
        \register[18][20] ), .D(\register[19][20] ), .S0(n1483), .S1(n1442), 
        .Y(n1296) );
  MXI4X1 U2237 ( .A(\register[0][21] ), .B(\register[1][21] ), .C(
        \register[2][21] ), .D(\register[3][21] ), .S0(n1484), .S1(n1443), .Y(
        n1308) );
  MXI4X1 U2238 ( .A(\register[16][21] ), .B(\register[17][21] ), .C(
        \register[18][21] ), .D(\register[19][21] ), .S0(n1483), .S1(n1442), 
        .Y(n1304) );
  MXI4X1 U2239 ( .A(\register[12][13] ), .B(\register[13][13] ), .C(
        \register[14][13] ), .D(\register[15][13] ), .S0(n1478), .S1(n1437), 
        .Y(n1241) );
  MXI4X1 U2240 ( .A(\register[12][14] ), .B(\register[13][14] ), .C(
        \register[14][14] ), .D(\register[15][14] ), .S0(n1479), .S1(n1438), 
        .Y(n1249) );
  MXI4X1 U2241 ( .A(\register[12][16] ), .B(\register[13][16] ), .C(
        \register[14][16] ), .D(\register[15][16] ), .S0(n1480), .S1(n1439), 
        .Y(n1265) );
  MXI4X1 U2242 ( .A(\register[12][15] ), .B(\register[13][15] ), .C(
        \register[14][15] ), .D(\register[15][15] ), .S0(n1480), .S1(n1439), 
        .Y(n1257) );
  MXI4X1 U2243 ( .A(\register[12][17] ), .B(\register[13][17] ), .C(
        \register[14][17] ), .D(\register[15][17] ), .S0(n1481), .S1(n1440), 
        .Y(n1273) );
  MXI4X1 U2244 ( .A(\register[12][18] ), .B(\register[13][18] ), .C(
        \register[14][18] ), .D(\register[15][18] ), .S0(n1482), .S1(n1441), 
        .Y(n1281) );
  MXI4X1 U2245 ( .A(\register[12][19] ), .B(\register[13][19] ), .C(
        \register[14][19] ), .D(\register[15][19] ), .S0(n1482), .S1(n1441), 
        .Y(n1289) );
  MXI4X1 U2246 ( .A(\register[12][20] ), .B(\register[13][20] ), .C(
        \register[14][20] ), .D(\register[15][20] ), .S0(n1483), .S1(n1442), 
        .Y(n1297) );
  MXI4X1 U2247 ( .A(\register[12][21] ), .B(\register[13][21] ), .C(
        \register[14][21] ), .D(\register[15][21] ), .S0(n1484), .S1(n1443), 
        .Y(n1305) );
  MXI4X1 U2248 ( .A(\register[8][13] ), .B(\register[9][13] ), .C(
        \register[10][13] ), .D(\register[11][13] ), .S0(n1478), .S1(n1437), 
        .Y(n1242) );
  MXI4X1 U2249 ( .A(\register[24][13] ), .B(\register[25][13] ), .C(
        \register[26][13] ), .D(\register[27][13] ), .S0(n1478), .S1(n1437), 
        .Y(n1238) );
  MXI4X1 U2250 ( .A(\register[8][14] ), .B(\register[9][14] ), .C(
        \register[10][14] ), .D(\register[11][14] ), .S0(n1479), .S1(n1438), 
        .Y(n1250) );
  MXI4X1 U2251 ( .A(\register[24][14] ), .B(\register[25][14] ), .C(
        \register[26][14] ), .D(\register[27][14] ), .S0(n1479), .S1(n1438), 
        .Y(n1246) );
  MXI4X1 U2252 ( .A(\register[8][16] ), .B(\register[9][16] ), .C(
        \register[10][16] ), .D(\register[11][16] ), .S0(n1480), .S1(n1439), 
        .Y(n1266) );
  MXI4X1 U2253 ( .A(\register[24][16] ), .B(\register[25][16] ), .C(
        \register[26][16] ), .D(\register[27][16] ), .S0(n1480), .S1(n1439), 
        .Y(n1262) );
  MXI4X1 U2254 ( .A(\register[8][15] ), .B(\register[9][15] ), .C(
        \register[10][15] ), .D(\register[11][15] ), .S0(n1480), .S1(n1439), 
        .Y(n1258) );
  MXI4X1 U2255 ( .A(\register[24][15] ), .B(\register[25][15] ), .C(
        \register[26][15] ), .D(\register[27][15] ), .S0(n1479), .S1(n1438), 
        .Y(n1254) );
  MXI4X1 U2256 ( .A(\register[8][17] ), .B(\register[9][17] ), .C(
        \register[10][17] ), .D(\register[11][17] ), .S0(n1481), .S1(n1440), 
        .Y(n1274) );
  MXI4X1 U2257 ( .A(\register[24][17] ), .B(\register[25][17] ), .C(
        \register[26][17] ), .D(\register[27][17] ), .S0(n1481), .S1(n1440), 
        .Y(n1270) );
  MXI4X1 U2258 ( .A(\register[8][18] ), .B(\register[9][18] ), .C(
        \register[10][18] ), .D(\register[11][18] ), .S0(n1482), .S1(n1441), 
        .Y(n1282) );
  MXI4X1 U2259 ( .A(\register[24][18] ), .B(\register[25][18] ), .C(
        \register[26][18] ), .D(\register[27][18] ), .S0(n1481), .S1(n1440), 
        .Y(n1278) );
  MXI4X1 U2260 ( .A(\register[8][19] ), .B(\register[9][19] ), .C(
        \register[10][19] ), .D(\register[11][19] ), .S0(n1482), .S1(n1441), 
        .Y(n1290) );
  MXI4X1 U2261 ( .A(\register[24][19] ), .B(\register[25][19] ), .C(
        \register[26][19] ), .D(\register[27][19] ), .S0(n1482), .S1(n1441), 
        .Y(n1286) );
  MXI4X1 U2262 ( .A(\register[8][20] ), .B(\register[9][20] ), .C(
        \register[10][20] ), .D(\register[11][20] ), .S0(n1483), .S1(n1442), 
        .Y(n1298) );
  MXI4X1 U2263 ( .A(\register[24][20] ), .B(\register[25][20] ), .C(
        \register[26][20] ), .D(\register[27][20] ), .S0(n1483), .S1(n1442), 
        .Y(n1294) );
  MXI4X1 U2264 ( .A(\register[8][21] ), .B(\register[9][21] ), .C(
        \register[10][21] ), .D(\register[11][21] ), .S0(n1484), .S1(n1443), 
        .Y(n1306) );
  MXI4X1 U2265 ( .A(\register[24][21] ), .B(\register[25][21] ), .C(
        \register[26][21] ), .D(\register[27][21] ), .S0(n1483), .S1(n1442), 
        .Y(n1302) );
  MX4X1 U2266 ( .A(n1312), .B(n1310), .C(n1311), .D(n1309), .S0(n1398), .S1(
        n1406), .Y(n1114) );
  MX4X1 U2267 ( .A(n1316), .B(n1314), .C(n1315), .D(n1313), .S0(n1398), .S1(
        n1406), .Y(n1113) );
  MXI4X1 U2268 ( .A(\register[28][22] ), .B(\register[29][22] ), .C(
        \register[30][22] ), .D(\register[31][22] ), .S0(n1484), .S1(n1443), 
        .Y(n1309) );
  MX4X1 U2269 ( .A(n1384), .B(n1382), .C(n1383), .D(n1381), .S0(n1399), .S1(
        n1407), .Y(n1132) );
  MX4X1 U2270 ( .A(n1388), .B(n1386), .C(n1387), .D(n1385), .S0(n1399), .S1(
        n1407), .Y(n1131) );
  MXI4X1 U2271 ( .A(\register[28][31] ), .B(\register[29][31] ), .C(
        \register[30][31] ), .D(\register[31][31] ), .S0(n1490), .S1(n1449), 
        .Y(n1381) );
  MX4X1 U2272 ( .A(n1332), .B(n1330), .C(n1331), .D(n1329), .S0(n1398), .S1(
        n1406), .Y(n1117) );
  MX4X1 U2273 ( .A(n1328), .B(n1326), .C(n1327), .D(n1325), .S0(n1398), .S1(
        n1406), .Y(n1118) );
  MXI4X1 U2274 ( .A(\register[0][24] ), .B(\register[1][24] ), .C(
        \register[2][24] ), .D(\register[3][24] ), .S0(n1486), .S1(n1445), .Y(
        n1332) );
  MX4X1 U2275 ( .A(n1340), .B(n1338), .C(n1339), .D(n1337), .S0(n1398), .S1(
        n1407), .Y(n1119) );
  MX4X1 U2276 ( .A(n1336), .B(n1334), .C(n1335), .D(n1333), .S0(n1398), .S1(
        n1406), .Y(n1120) );
  MXI4X1 U2277 ( .A(\register[0][25] ), .B(\register[1][25] ), .C(
        \register[2][25] ), .D(\register[3][25] ), .S0(n1486), .S1(n1445), .Y(
        n1340) );
  MX4X1 U2278 ( .A(n1380), .B(n1378), .C(n1379), .D(n1377), .S0(n1399), .S1(
        n1407), .Y(n1129) );
  MX4X1 U2279 ( .A(n1376), .B(n1374), .C(n1375), .D(n1373), .S0(n1399), .S1(
        n1407), .Y(n1130) );
  MXI4X1 U2280 ( .A(\register[0][30] ), .B(\register[1][30] ), .C(
        \register[2][30] ), .D(\register[3][30] ), .S0(n1490), .S1(n1449), .Y(
        n1380) );
  MX4X1 U2281 ( .A(n1368), .B(n1366), .C(n1367), .D(n1365), .S0(n1399), .S1(
        n1407), .Y(n1128) );
  MX4X1 U2282 ( .A(n1372), .B(n1370), .C(n1371), .D(n1369), .S0(n1399), .S1(
        n1407), .Y(n1127) );
  MXI4X1 U2283 ( .A(\register[28][29] ), .B(\register[29][29] ), .C(
        \register[30][29] ), .D(\register[31][29] ), .S0(n1489), .S1(n1448), 
        .Y(n1365) );
  MX4X1 U2284 ( .A(n1320), .B(n1318), .C(n1319), .D(n1317), .S0(n1398), .S1(
        n1406), .Y(n1116) );
  MX4X1 U2285 ( .A(n1324), .B(n1322), .C(n1323), .D(n1321), .S0(n1398), .S1(
        n1406), .Y(n1115) );
  MXI4X1 U2286 ( .A(\register[28][23] ), .B(\register[29][23] ), .C(
        \register[30][23] ), .D(\register[31][23] ), .S0(n1485), .S1(n1444), 
        .Y(n1317) );
  MX4X1 U2287 ( .A(n1344), .B(n1342), .C(n1343), .D(n1341), .S0(n1399), .S1(
        n1407), .Y(n1122) );
  MX4X1 U2288 ( .A(n1348), .B(n1346), .C(n1347), .D(n1345), .S0(n1399), .S1(
        n1407), .Y(n1121) );
  MXI4X1 U2289 ( .A(\register[28][26] ), .B(\register[29][26] ), .C(
        \register[30][26] ), .D(\register[31][26] ), .S0(n1487), .S1(n1446), 
        .Y(n1341) );
  MX4X1 U2290 ( .A(n1356), .B(n1354), .C(n1355), .D(n1353), .S0(n1399), .S1(
        n1407), .Y(n1123) );
  MX4X1 U2291 ( .A(n1352), .B(n1350), .C(n1351), .D(n1349), .S0(n1399), .S1(
        n1407), .Y(n1124) );
  MXI4X1 U2292 ( .A(\register[8][27] ), .B(\register[9][27] ), .C(
        \register[10][27] ), .D(\register[11][27] ), .S0(n1488), .S1(n1447), 
        .Y(n1354) );
  MX4X1 U2293 ( .A(n1364), .B(n1362), .C(n1363), .D(n1361), .S0(n1399), .S1(
        n1407), .Y(n1125) );
  MX4X1 U2294 ( .A(n1360), .B(n1358), .C(n1359), .D(n1357), .S0(n1399), .S1(
        n1407), .Y(n1126) );
  MXI4X1 U2295 ( .A(\register[0][28] ), .B(\register[1][28] ), .C(
        \register[2][28] ), .D(\register[3][28] ), .S0(n1488), .S1(n1447), .Y(
        n1364) );
  MXI4X1 U2296 ( .A(\register[4][22] ), .B(\register[5][22] ), .C(
        \register[6][22] ), .D(\register[7][22] ), .S0(n1484), .S1(n1443), .Y(
        n1315) );
  MXI4X1 U2297 ( .A(\register[20][22] ), .B(\register[21][22] ), .C(
        \register[22][22] ), .D(\register[23][22] ), .S0(n1484), .S1(n1443), 
        .Y(n1311) );
  MXI4X1 U2298 ( .A(\register[4][23] ), .B(\register[5][23] ), .C(
        \register[6][23] ), .D(\register[7][23] ), .S0(n1485), .S1(n1444), .Y(
        n1323) );
  MXI4X1 U2299 ( .A(\register[20][23] ), .B(\register[21][23] ), .C(
        \register[22][23] ), .D(\register[23][23] ), .S0(n1485), .S1(n1444), 
        .Y(n1319) );
  MXI4X1 U2300 ( .A(\register[20][24] ), .B(\register[21][24] ), .C(
        \register[22][24] ), .D(\register[23][24] ), .S0(n1485), .S1(n1444), 
        .Y(n1327) );
  MXI4X1 U2301 ( .A(\register[4][24] ), .B(\register[5][24] ), .C(
        \register[6][24] ), .D(\register[7][24] ), .S0(n1486), .S1(n1445), .Y(
        n1331) );
  MXI4X1 U2302 ( .A(\register[20][25] ), .B(\register[21][25] ), .C(
        \register[22][25] ), .D(\register[23][25] ), .S0(n1486), .S1(n1445), 
        .Y(n1335) );
  MXI4X1 U2303 ( .A(\register[4][25] ), .B(\register[5][25] ), .C(
        \register[6][25] ), .D(\register[7][25] ), .S0(n1486), .S1(n1445), .Y(
        n1339) );
  MXI4X1 U2304 ( .A(\register[4][26] ), .B(\register[5][26] ), .C(
        \register[6][26] ), .D(\register[7][26] ), .S0(n1487), .S1(n1446), .Y(
        n1347) );
  MXI4X1 U2305 ( .A(\register[20][26] ), .B(\register[21][26] ), .C(
        \register[22][26] ), .D(\register[23][26] ), .S0(n1487), .S1(n1446), 
        .Y(n1343) );
  MXI4X1 U2306 ( .A(\register[20][27] ), .B(\register[21][27] ), .C(
        \register[22][27] ), .D(\register[23][27] ), .S0(n1487), .S1(n1446), 
        .Y(n1351) );
  MXI4X1 U2307 ( .A(\register[4][27] ), .B(\register[5][27] ), .C(
        \register[6][27] ), .D(\register[7][27] ), .S0(n1488), .S1(n1447), .Y(
        n1355) );
  MXI4X1 U2308 ( .A(\register[20][30] ), .B(\register[21][30] ), .C(
        \register[22][30] ), .D(\register[23][30] ), .S0(n1489), .S1(n1448), 
        .Y(n1375) );
  MXI4X1 U2309 ( .A(\register[4][30] ), .B(\register[5][30] ), .C(
        \register[6][30] ), .D(\register[7][30] ), .S0(n1490), .S1(n1449), .Y(
        n1379) );
  MXI4X1 U2310 ( .A(\register[20][28] ), .B(\register[21][28] ), .C(
        \register[22][28] ), .D(\register[23][28] ), .S0(n1488), .S1(n1447), 
        .Y(n1359) );
  MXI4X1 U2311 ( .A(\register[4][28] ), .B(\register[5][28] ), .C(
        \register[6][28] ), .D(\register[7][28] ), .S0(n1488), .S1(n1447), .Y(
        n1363) );
  MXI4X1 U2312 ( .A(\register[4][29] ), .B(\register[5][29] ), .C(
        \register[6][29] ), .D(\register[7][29] ), .S0(n1489), .S1(n1448), .Y(
        n1371) );
  MXI4X1 U2313 ( .A(\register[20][29] ), .B(\register[21][29] ), .C(
        \register[22][29] ), .D(\register[23][29] ), .S0(n1489), .S1(n1448), 
        .Y(n1367) );
  MXI4X1 U2314 ( .A(\register[4][31] ), .B(\register[5][31] ), .C(
        \register[6][31] ), .D(\register[7][31] ), .S0(n1490), .S1(n1449), .Y(
        n1387) );
  MXI4X1 U2315 ( .A(\register[20][31] ), .B(\register[21][31] ), .C(
        \register[22][31] ), .D(\register[23][31] ), .S0(n1490), .S1(n1449), 
        .Y(n1383) );
  MXI4X1 U2316 ( .A(\register[0][22] ), .B(\register[1][22] ), .C(
        \register[2][22] ), .D(\register[3][22] ), .S0(n1484), .S1(n1443), .Y(
        n1316) );
  MXI4X1 U2317 ( .A(\register[16][22] ), .B(\register[17][22] ), .C(
        \register[18][22] ), .D(\register[19][22] ), .S0(n1484), .S1(n1443), 
        .Y(n1312) );
  MXI4X1 U2318 ( .A(\register[0][23] ), .B(\register[1][23] ), .C(
        \register[2][23] ), .D(\register[3][23] ), .S0(n1485), .S1(n1444), .Y(
        n1324) );
  MXI4X1 U2319 ( .A(\register[16][23] ), .B(\register[17][23] ), .C(
        \register[18][23] ), .D(\register[19][23] ), .S0(n1485), .S1(n1444), 
        .Y(n1320) );
  MXI4X1 U2320 ( .A(\register[16][24] ), .B(\register[17][24] ), .C(
        \register[18][24] ), .D(\register[19][24] ), .S0(n1485), .S1(n1444), 
        .Y(n1328) );
  MXI4X1 U2321 ( .A(\register[16][25] ), .B(\register[17][25] ), .C(
        \register[18][25] ), .D(\register[19][25] ), .S0(n1486), .S1(n1445), 
        .Y(n1336) );
  MXI4X1 U2322 ( .A(\register[0][26] ), .B(\register[1][26] ), .C(
        \register[2][26] ), .D(\register[3][26] ), .S0(n1487), .S1(n1446), .Y(
        n1348) );
  MXI4X1 U2323 ( .A(\register[16][26] ), .B(\register[17][26] ), .C(
        \register[18][26] ), .D(\register[19][26] ), .S0(n1487), .S1(n1446), 
        .Y(n1344) );
  MXI4X1 U2324 ( .A(\register[16][27] ), .B(\register[17][27] ), .C(
        \register[18][27] ), .D(\register[19][27] ), .S0(n1487), .S1(n1446), 
        .Y(n1352) );
  MXI4X1 U2325 ( .A(\register[0][27] ), .B(\register[1][27] ), .C(
        \register[2][27] ), .D(\register[3][27] ), .S0(n1488), .S1(n1447), .Y(
        n1356) );
  MXI4X1 U2326 ( .A(\register[16][30] ), .B(\register[17][30] ), .C(
        \register[18][30] ), .D(\register[19][30] ), .S0(n1489), .S1(n1448), 
        .Y(n1376) );
  MXI4X1 U2327 ( .A(\register[16][28] ), .B(\register[17][28] ), .C(
        \register[18][28] ), .D(\register[19][28] ), .S0(n1488), .S1(n1447), 
        .Y(n1360) );
  MXI4X1 U2328 ( .A(\register[0][29] ), .B(\register[1][29] ), .C(
        \register[2][29] ), .D(\register[3][29] ), .S0(n1489), .S1(n1448), .Y(
        n1372) );
  MXI4X1 U2329 ( .A(\register[16][29] ), .B(\register[17][29] ), .C(
        \register[18][29] ), .D(\register[19][29] ), .S0(n1489), .S1(n1448), 
        .Y(n1368) );
  MXI4X1 U2330 ( .A(\register[0][31] ), .B(\register[1][31] ), .C(
        \register[2][31] ), .D(\register[3][31] ), .S0(n1490), .S1(n1449), .Y(
        n1388) );
  MXI4X1 U2331 ( .A(\register[16][31] ), .B(\register[17][31] ), .C(
        \register[18][31] ), .D(\register[19][31] ), .S0(n1490), .S1(n1449), 
        .Y(n1384) );
  MXI4X1 U2332 ( .A(\register[12][22] ), .B(\register[13][22] ), .C(
        \register[14][22] ), .D(\register[15][22] ), .S0(n1484), .S1(n1443), 
        .Y(n1313) );
  MXI4X1 U2333 ( .A(\register[12][23] ), .B(\register[13][23] ), .C(
        \register[14][23] ), .D(\register[15][23] ), .S0(n1485), .S1(n1444), 
        .Y(n1321) );
  MXI4X1 U2334 ( .A(\register[28][24] ), .B(\register[29][24] ), .C(
        \register[30][24] ), .D(\register[31][24] ), .S0(n1485), .S1(n1444), 
        .Y(n1325) );
  MXI4X1 U2335 ( .A(\register[12][24] ), .B(\register[13][24] ), .C(
        \register[14][24] ), .D(\register[15][24] ), .S0(n1486), .S1(n1445), 
        .Y(n1329) );
  MXI4X1 U2336 ( .A(\register[28][25] ), .B(\register[29][25] ), .C(
        \register[30][25] ), .D(\register[31][25] ), .S0(n1486), .S1(n1445), 
        .Y(n1333) );
  MXI4X1 U2337 ( .A(\register[12][25] ), .B(\register[13][25] ), .C(
        \register[14][25] ), .D(\register[15][25] ), .S0(n1486), .S1(n1445), 
        .Y(n1337) );
  MXI4X1 U2338 ( .A(\register[12][26] ), .B(\register[13][26] ), .C(
        \register[14][26] ), .D(\register[15][26] ), .S0(n1487), .S1(n1446), 
        .Y(n1345) );
  MXI4X1 U2339 ( .A(\register[28][27] ), .B(\register[29][27] ), .C(
        \register[30][27] ), .D(\register[31][27] ), .S0(n1487), .S1(n1446), 
        .Y(n1349) );
  MXI4X1 U2340 ( .A(\register[12][27] ), .B(\register[13][27] ), .C(
        \register[14][27] ), .D(\register[15][27] ), .S0(n1488), .S1(n1447), 
        .Y(n1353) );
  MXI4X1 U2341 ( .A(\register[28][30] ), .B(\register[29][30] ), .C(
        \register[30][30] ), .D(\register[31][30] ), .S0(n1489), .S1(n1448), 
        .Y(n1373) );
  MXI4X1 U2342 ( .A(\register[12][30] ), .B(\register[13][30] ), .C(
        \register[14][30] ), .D(\register[15][30] ), .S0(n1490), .S1(n1449), 
        .Y(n1377) );
  MXI4X1 U2343 ( .A(\register[28][28] ), .B(\register[29][28] ), .C(
        \register[30][28] ), .D(\register[31][28] ), .S0(n1488), .S1(n1447), 
        .Y(n1357) );
  MXI4X1 U2344 ( .A(\register[12][28] ), .B(\register[13][28] ), .C(
        \register[14][28] ), .D(\register[15][28] ), .S0(n1488), .S1(n1447), 
        .Y(n1361) );
  MXI4X1 U2345 ( .A(\register[12][29] ), .B(\register[13][29] ), .C(
        \register[14][29] ), .D(\register[15][29] ), .S0(n1489), .S1(n1448), 
        .Y(n1369) );
  MXI4X1 U2346 ( .A(\register[12][31] ), .B(\register[13][31] ), .C(
        \register[14][31] ), .D(\register[15][31] ), .S0(n1490), .S1(n1449), 
        .Y(n1385) );
  MXI4X1 U2347 ( .A(\register[8][22] ), .B(\register[9][22] ), .C(
        \register[10][22] ), .D(\register[11][22] ), .S0(n1484), .S1(n1443), 
        .Y(n1314) );
  MXI4X1 U2348 ( .A(\register[24][22] ), .B(\register[25][22] ), .C(
        \register[26][22] ), .D(\register[27][22] ), .S0(n1484), .S1(n1443), 
        .Y(n1310) );
  MXI4X1 U2349 ( .A(\register[8][23] ), .B(\register[9][23] ), .C(
        \register[10][23] ), .D(\register[11][23] ), .S0(n1485), .S1(n1444), 
        .Y(n1322) );
  MXI4X1 U2350 ( .A(\register[24][23] ), .B(\register[25][23] ), .C(
        \register[26][23] ), .D(\register[27][23] ), .S0(n1485), .S1(n1444), 
        .Y(n1318) );
  MXI4X1 U2351 ( .A(\register[24][24] ), .B(\register[25][24] ), .C(
        \register[26][24] ), .D(\register[27][24] ), .S0(n1485), .S1(n1444), 
        .Y(n1326) );
  MXI4X1 U2352 ( .A(\register[8][24] ), .B(\register[9][24] ), .C(
        \register[10][24] ), .D(\register[11][24] ), .S0(n1486), .S1(n1445), 
        .Y(n1330) );
  MXI4X1 U2353 ( .A(\register[24][25] ), .B(\register[25][25] ), .C(
        \register[26][25] ), .D(\register[27][25] ), .S0(n1486), .S1(n1445), 
        .Y(n1334) );
  MXI4X1 U2354 ( .A(\register[8][25] ), .B(\register[9][25] ), .C(
        \register[10][25] ), .D(\register[11][25] ), .S0(n1486), .S1(n1445), 
        .Y(n1338) );
  MXI4X1 U2355 ( .A(\register[8][26] ), .B(\register[9][26] ), .C(
        \register[10][26] ), .D(\register[11][26] ), .S0(n1487), .S1(n1446), 
        .Y(n1346) );
  MXI4X1 U2356 ( .A(\register[24][26] ), .B(\register[25][26] ), .C(
        \register[26][26] ), .D(\register[27][26] ), .S0(n1487), .S1(n1446), 
        .Y(n1342) );
  MXI4X1 U2357 ( .A(\register[24][27] ), .B(\register[25][27] ), .C(
        \register[26][27] ), .D(\register[27][27] ), .S0(n1487), .S1(n1446), 
        .Y(n1350) );
  MXI4X1 U2358 ( .A(\register[24][30] ), .B(\register[25][30] ), .C(
        \register[26][30] ), .D(\register[27][30] ), .S0(n1489), .S1(n1448), 
        .Y(n1374) );
  MXI4X1 U2359 ( .A(\register[8][30] ), .B(\register[9][30] ), .C(
        \register[10][30] ), .D(\register[11][30] ), .S0(n1490), .S1(n1449), 
        .Y(n1378) );
  MXI4X1 U2360 ( .A(\register[24][28] ), .B(\register[25][28] ), .C(
        \register[26][28] ), .D(\register[27][28] ), .S0(n1488), .S1(n1447), 
        .Y(n1358) );
  MXI4X1 U2361 ( .A(\register[8][28] ), .B(\register[9][28] ), .C(
        \register[10][28] ), .D(\register[11][28] ), .S0(n1488), .S1(n1447), 
        .Y(n1362) );
  MXI4X1 U2362 ( .A(\register[8][29] ), .B(\register[9][29] ), .C(
        \register[10][29] ), .D(\register[11][29] ), .S0(n1489), .S1(n1448), 
        .Y(n1370) );
  MXI4X1 U2363 ( .A(\register[24][29] ), .B(\register[25][29] ), .C(
        \register[26][29] ), .D(\register[27][29] ), .S0(n1489), .S1(n1448), 
        .Y(n1366) );
  MXI4X1 U2364 ( .A(\register[8][31] ), .B(\register[9][31] ), .C(
        \register[10][31] ), .D(\register[11][31] ), .S0(n1490), .S1(n1449), 
        .Y(n1386) );
  MXI4X1 U2365 ( .A(\register[24][31] ), .B(\register[25][31] ), .C(
        \register[26][31] ), .D(\register[27][31] ), .S0(n1490), .S1(n1449), 
        .Y(n1382) );
  CLKBUFX3 U2366 ( .A(n1392), .Y(n1389) );
  CLKBUFX3 U2367 ( .A(N14), .Y(n1392) );
  CLKBUFX3 U2368 ( .A(n1816), .Y(n1813) );
  CLKBUFX3 U2369 ( .A(N19), .Y(n1816) );
  CLKBUFX3 U2370 ( .A(n1408), .Y(n1403) );
  CLKBUFX3 U2371 ( .A(N12), .Y(n1408) );
  CLKBUFX3 U2372 ( .A(N14), .Y(n1393) );
  CLKBUFX3 U2373 ( .A(N12), .Y(n1409) );
  CLKBUFX3 U2374 ( .A(N12), .Y(n1410) );
  CLKBUFX3 U2375 ( .A(N19), .Y(n1817) );
endmodule


module Mux_WIDTH5_0 ( data1_i, data2_i, select_i, data_o );
  input [4:0] data1_i;
  input [4:0] data2_i;
  output [4:0] data_o;
  input select_i;
  wire   n1;

  CLKINVX1 U1 ( .A(select_i), .Y(n1) );
  AO22X1 U2 ( .A0(data2_i[1]), .A1(select_i), .B0(data1_i[1]), .B1(n1), .Y(
        data_o[1]) );
  AO22X1 U3 ( .A0(data2_i[0]), .A1(select_i), .B0(data1_i[0]), .B1(n1), .Y(
        data_o[0]) );
  AO22X1 U4 ( .A0(data2_i[2]), .A1(select_i), .B0(data1_i[2]), .B1(n1), .Y(
        data_o[2]) );
  AO22X1 U5 ( .A0(select_i), .A1(data2_i[4]), .B0(data1_i[4]), .B1(n1), .Y(
        data_o[4]) );
  AO22X1 U6 ( .A0(data2_i[3]), .A1(select_i), .B0(data1_i[3]), .B1(n1), .Y(
        data_o[3]) );
endmodule


module Mux_WIDTH32_0 ( data1_i, data2_i, select_i, data_o );
  input [31:0] data1_i;
  input [31:0] data2_i;
  output [31:0] data_o;
  input select_i;
  wire   n1, n2, n3, n4, n5, n6, n7;

  AO22X1 U1 ( .A0(data2_i[19]), .A1(select_i), .B0(data1_i[19]), .B1(n5), .Y(
        data_o[19]) );
  AO22X1 U2 ( .A0(data2_i[20]), .A1(select_i), .B0(data1_i[20]), .B1(n5), .Y(
        data_o[20]) );
  AO22X1 U3 ( .A0(data2_i[21]), .A1(n1), .B0(data1_i[21]), .B1(n5), .Y(
        data_o[21]) );
  AO22X1 U4 ( .A0(data2_i[26]), .A1(select_i), .B0(data1_i[26]), .B1(n5), .Y(
        data_o[26]) );
  AO22X1 U5 ( .A0(data2_i[27]), .A1(n1), .B0(data1_i[27]), .B1(n5), .Y(
        data_o[27]) );
  AO22X1 U6 ( .A0(data2_i[28]), .A1(select_i), .B0(data1_i[28]), .B1(n5), .Y(
        data_o[28]) );
  AO22X1 U7 ( .A0(data2_i[29]), .A1(n1), .B0(data1_i[29]), .B1(n5), .Y(
        data_o[29]) );
  CLKBUFX3 U8 ( .A(n7), .Y(n4) );
  CLKBUFX3 U9 ( .A(n4), .Y(n2) );
  CLKBUFX3 U10 ( .A(n7), .Y(n3) );
  CLKBUFX3 U11 ( .A(n7), .Y(n5) );
  CLKBUFX3 U12 ( .A(n7), .Y(n6) );
  CLKINVX1 U13 ( .A(n1), .Y(n7) );
  AO22X1 U14 ( .A0(data2_i[1]), .A1(n1), .B0(data1_i[1]), .B1(n5), .Y(
        data_o[1]) );
  AO22X1 U15 ( .A0(data2_i[2]), .A1(select_i), .B0(data1_i[2]), .B1(n5), .Y(
        data_o[2]) );
  AO22X1 U16 ( .A0(data2_i[3]), .A1(n1), .B0(data1_i[3]), .B1(n6), .Y(
        data_o[3]) );
  AO22X1 U17 ( .A0(data2_i[0]), .A1(select_i), .B0(data1_i[0]), .B1(n2), .Y(
        data_o[0]) );
  AO22X1 U18 ( .A0(data2_i[8]), .A1(select_i), .B0(data1_i[8]), .B1(n6), .Y(
        data_o[8]) );
  AO22X1 U19 ( .A0(data2_i[4]), .A1(n1), .B0(data1_i[4]), .B1(n6), .Y(
        data_o[4]) );
  AO22X1 U20 ( .A0(data2_i[5]), .A1(select_i), .B0(data1_i[5]), .B1(n6), .Y(
        data_o[5]) );
  AO22X1 U21 ( .A0(data2_i[6]), .A1(n1), .B0(data1_i[6]), .B1(n6), .Y(
        data_o[6]) );
  AO22X1 U22 ( .A0(data2_i[7]), .A1(select_i), .B0(data1_i[7]), .B1(n6), .Y(
        data_o[7]) );
  AO22X1 U23 ( .A0(select_i), .A1(data2_i[9]), .B0(data1_i[9]), .B1(n6), .Y(
        data_o[9]) );
  AO22X1 U24 ( .A0(data2_i[10]), .A1(n1), .B0(data1_i[10]), .B1(n2), .Y(
        data_o[10]) );
  AO22X1 U25 ( .A0(data2_i[11]), .A1(select_i), .B0(data1_i[11]), .B1(n3), .Y(
        data_o[11]) );
  AO22X1 U26 ( .A0(data2_i[12]), .A1(n1), .B0(data1_i[12]), .B1(n3), .Y(
        data_o[12]) );
  AO22X1 U27 ( .A0(data2_i[13]), .A1(select_i), .B0(data1_i[13]), .B1(n4), .Y(
        data_o[13]) );
  AO22X1 U28 ( .A0(data2_i[18]), .A1(n1), .B0(data1_i[18]), .B1(n5), .Y(
        data_o[18]) );
  AO22X1 U29 ( .A0(data2_i[15]), .A1(select_i), .B0(data1_i[15]), .B1(n5), .Y(
        data_o[15]) );
  AO22X1 U30 ( .A0(data2_i[16]), .A1(n1), .B0(data1_i[16]), .B1(n5), .Y(
        data_o[16]) );
  AO22X1 U31 ( .A0(data2_i[17]), .A1(select_i), .B0(data1_i[17]), .B1(n5), .Y(
        data_o[17]) );
  AO22X1 U32 ( .A0(data2_i[22]), .A1(n1), .B0(data1_i[22]), .B1(n5), .Y(
        data_o[22]) );
  AO22X1 U33 ( .A0(data2_i[14]), .A1(n1), .B0(data1_i[14]), .B1(n4), .Y(
        data_o[14]) );
  AO22X1 U34 ( .A0(data2_i[23]), .A1(select_i), .B0(data1_i[23]), .B1(n5), .Y(
        data_o[23]) );
  AO22X1 U35 ( .A0(data2_i[24]), .A1(n1), .B0(data1_i[24]), .B1(n5), .Y(
        data_o[24]) );
  AO22X1 U36 ( .A0(data2_i[25]), .A1(select_i), .B0(data1_i[25]), .B1(n5), .Y(
        data_o[25]) );
  AO22X1 U37 ( .A0(data2_i[30]), .A1(n1), .B0(data1_i[30]), .B1(n6), .Y(
        data_o[30]) );
  AO22X1 U38 ( .A0(data2_i[31]), .A1(n1), .B0(data1_i[31]), .B1(n6), .Y(
        data_o[31]) );
  CLKBUFX3 U39 ( .A(select_i), .Y(n1) );
endmodule


module Mux_WIDTH32_5 ( data1_i, data2_i, select_i, data_o );
  input [31:0] data1_i;
  input [31:0] data2_i;
  output [31:0] data_o;
  input select_i;
  wire   n1, n2, n3, n4, n5, n6, n7;

  CLKBUFX3 U1 ( .A(n7), .Y(n4) );
  CLKBUFX3 U2 ( .A(n4), .Y(n2) );
  CLKBUFX3 U3 ( .A(n7), .Y(n3) );
  CLKBUFX3 U4 ( .A(n7), .Y(n5) );
  CLKBUFX3 U5 ( .A(n7), .Y(n6) );
  CLKINVX1 U6 ( .A(n1), .Y(n7) );
  CLKBUFX3 U7 ( .A(select_i), .Y(n1) );
  AO22X1 U8 ( .A0(data2_i[1]), .A1(select_i), .B0(data1_i[1]), .B1(n5), .Y(
        data_o[1]) );
  AO22X1 U9 ( .A0(data2_i[2]), .A1(select_i), .B0(data1_i[2]), .B1(n5), .Y(
        data_o[2]) );
  AO22X1 U10 ( .A0(data2_i[15]), .A1(n1), .B0(data1_i[15]), .B1(n5), .Y(
        data_o[15]) );
  AO22X1 U11 ( .A0(data2_i[16]), .A1(select_i), .B0(data1_i[16]), .B1(n5), .Y(
        data_o[16]) );
  AO22X1 U12 ( .A0(data2_i[17]), .A1(n1), .B0(data1_i[17]), .B1(n5), .Y(
        data_o[17]) );
  AO22X1 U13 ( .A0(data2_i[18]), .A1(select_i), .B0(data1_i[18]), .B1(n5), .Y(
        data_o[18]) );
  AO22X1 U14 ( .A0(data2_i[19]), .A1(n1), .B0(data1_i[19]), .B1(n5), .Y(
        data_o[19]) );
  AO22X1 U15 ( .A0(data2_i[20]), .A1(n1), .B0(data1_i[20]), .B1(n5), .Y(
        data_o[20]) );
  AO22X1 U16 ( .A0(data2_i[21]), .A1(select_i), .B0(data1_i[21]), .B1(n5), .Y(
        data_o[21]) );
  AO22X1 U17 ( .A0(data2_i[22]), .A1(n1), .B0(data1_i[22]), .B1(n5), .Y(
        data_o[22]) );
  AO22X1 U18 ( .A0(data2_i[23]), .A1(select_i), .B0(data1_i[23]), .B1(n5), .Y(
        data_o[23]) );
  AO22X1 U19 ( .A0(data2_i[24]), .A1(n1), .B0(data1_i[24]), .B1(n5), .Y(
        data_o[24]) );
  AO22X1 U20 ( .A0(data2_i[25]), .A1(select_i), .B0(data1_i[25]), .B1(n5), .Y(
        data_o[25]) );
  AO22X1 U21 ( .A0(data2_i[26]), .A1(n1), .B0(data1_i[26]), .B1(n5), .Y(
        data_o[26]) );
  AO22X1 U22 ( .A0(data2_i[27]), .A1(select_i), .B0(data1_i[27]), .B1(n5), .Y(
        data_o[27]) );
  AO22X1 U23 ( .A0(data2_i[28]), .A1(n1), .B0(data1_i[28]), .B1(n5), .Y(
        data_o[28]) );
  AO22X1 U24 ( .A0(data2_i[29]), .A1(select_i), .B0(data1_i[29]), .B1(n5), .Y(
        data_o[29]) );
  AO22X1 U25 ( .A0(data2_i[10]), .A1(select_i), .B0(data1_i[10]), .B1(n2), .Y(
        data_o[10]) );
  AO22X1 U26 ( .A0(data2_i[11]), .A1(n1), .B0(data1_i[11]), .B1(n3), .Y(
        data_o[11]) );
  AO22X1 U27 ( .A0(data2_i[12]), .A1(select_i), .B0(data1_i[12]), .B1(n3), .Y(
        data_o[12]) );
  AO22X1 U28 ( .A0(data2_i[13]), .A1(n1), .B0(data1_i[13]), .B1(n4), .Y(
        data_o[13]) );
  AO22X1 U29 ( .A0(data2_i[14]), .A1(select_i), .B0(data1_i[14]), .B1(n4), .Y(
        data_o[14]) );
  AO22X1 U30 ( .A0(data2_i[0]), .A1(n1), .B0(data1_i[0]), .B1(n2), .Y(
        data_o[0]) );
  AO22X1 U31 ( .A0(data2_i[3]), .A1(n1), .B0(data1_i[3]), .B1(n6), .Y(
        data_o[3]) );
  AO22X1 U32 ( .A0(data2_i[4]), .A1(select_i), .B0(data1_i[4]), .B1(n6), .Y(
        data_o[4]) );
  AO22X1 U33 ( .A0(data2_i[5]), .A1(n1), .B0(data1_i[5]), .B1(n6), .Y(
        data_o[5]) );
  AO22X1 U34 ( .A0(data2_i[6]), .A1(select_i), .B0(data1_i[6]), .B1(n6), .Y(
        data_o[6]) );
  AO22X1 U35 ( .A0(data2_i[7]), .A1(n1), .B0(data1_i[7]), .B1(n6), .Y(
        data_o[7]) );
  AO22X1 U36 ( .A0(data2_i[8]), .A1(select_i), .B0(data1_i[8]), .B1(n6), .Y(
        data_o[8]) );
  AO22X1 U37 ( .A0(n1), .A1(data2_i[9]), .B0(data1_i[9]), .B1(n6), .Y(
        data_o[9]) );
  AO22X1 U38 ( .A0(data2_i[30]), .A1(n1), .B0(data1_i[30]), .B1(n6), .Y(
        data_o[30]) );
  AO22X1 U39 ( .A0(data2_i[31]), .A1(n1), .B0(data1_i[31]), .B1(n6), .Y(
        data_o[31]) );
endmodule


module Add_ALU_0_DW01_add_0 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [31:1] carry;

  ADDFXL U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFXL U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFXL U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFXL U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFXL U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFXL U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFXL U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFXL U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFXL U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFXL U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFXL U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFXL U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFXL U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFXL U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFXL U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFXL U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFXL U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFXL U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFXL U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFXL U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFXL U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFXL U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFXL U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFXL U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFXL U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFXL U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFXL U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXL U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXL U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  XOR3X1 U1_31 ( .A(A[31]), .B(B[31]), .C(carry[31]), .Y(SUM[31]) );
  ADDFXL U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module Add_ALU_0 ( data1_i, data2_i, Add_ALU_o );
  input [31:0] data1_i;
  input [31:0] data2_i;
  output [31:0] Add_ALU_o;


  Add_ALU_0_DW01_add_0 add_269 ( .A(data1_i), .B(data2_i), .CI(1'b0), .SUM(
        Add_ALU_o) );
endmodule


module Add_ALU_1_DW01_add_0 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1, n2;
  wire   [31:1] carry;

  ADDFXL U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  XOR3X1 U1_31 ( .A(A[31]), .B(B[31]), .C(carry[31]), .Y(SUM[31]) );
  ADDFXL U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFXL U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  ADDFXL U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFXL U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFXL U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFXL U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFXL U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFXL U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFXL U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFXL U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFXL U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFXL U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFXL U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFXL U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFXL U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFXL U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFXL U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFXL U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFXL U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFXL U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFXL U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFXL U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFXL U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFXL U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFXL U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFXL U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFXL U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXL U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXL U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  CLKINVX1 U2 ( .A(A[0]), .Y(n2) );
  XNOR2X1 U3 ( .A(B[0]), .B(n2), .Y(SUM[0]) );
endmodule


module Add_ALU_1 ( data1_i, data2_i, Add_ALU_o );
  input [31:0] data1_i;
  input [31:0] data2_i;
  output [31:0] Add_ALU_o;


  Add_ALU_1_DW01_add_0 add_269 ( .A(data1_i), .B(data2_i), .CI(1'b0), .SUM(
        Add_ALU_o) );
endmodule


module Mux_WIDTH32_4 ( data1_i, data2_i, select_i, data_o );
  input [31:0] data1_i;
  input [31:0] data2_i;
  output [31:0] data_o;
  input select_i;
  wire   n1, n2, n3, n4, n5, n6, n7;

  CLKBUFX3 U1 ( .A(n7), .Y(n4) );
  CLKBUFX3 U2 ( .A(n7), .Y(n2) );
  CLKBUFX3 U3 ( .A(n7), .Y(n3) );
  CLKBUFX3 U4 ( .A(n7), .Y(n5) );
  CLKBUFX3 U5 ( .A(n7), .Y(n6) );
  CLKINVX1 U6 ( .A(n1), .Y(n7) );
  CLKBUFX3 U7 ( .A(select_i), .Y(n1) );
  AO22X1 U8 ( .A0(data2_i[31]), .A1(select_i), .B0(data1_i[31]), .B1(n6), .Y(
        data_o[31]) );
  AO22X1 U9 ( .A0(data2_i[30]), .A1(select_i), .B0(data1_i[30]), .B1(n6), .Y(
        data_o[30]) );
  AO22X1 U10 ( .A0(data2_i[18]), .A1(select_i), .B0(data1_i[18]), .B1(n5), .Y(
        data_o[18]) );
  AO22X1 U11 ( .A0(data2_i[19]), .A1(select_i), .B0(data1_i[19]), .B1(n5), .Y(
        data_o[19]) );
  AO22X1 U12 ( .A0(data2_i[20]), .A1(n1), .B0(data1_i[20]), .B1(n5), .Y(
        data_o[20]) );
  AO22X1 U13 ( .A0(data2_i[21]), .A1(select_i), .B0(data1_i[21]), .B1(n5), .Y(
        data_o[21]) );
  AO22X1 U14 ( .A0(data2_i[23]), .A1(select_i), .B0(data1_i[23]), .B1(n5), .Y(
        data_o[23]) );
  AO22X1 U15 ( .A0(data2_i[24]), .A1(select_i), .B0(data1_i[24]), .B1(n5), .Y(
        data_o[24]) );
  AO22X1 U16 ( .A0(data2_i[26]), .A1(select_i), .B0(data1_i[26]), .B1(n5), .Y(
        data_o[26]) );
  AO22X1 U17 ( .A0(data2_i[28]), .A1(select_i), .B0(data1_i[28]), .B1(n5), .Y(
        data_o[28]) );
  AO22X1 U18 ( .A0(data2_i[29]), .A1(select_i), .B0(data1_i[29]), .B1(n5), .Y(
        data_o[29]) );
  AO22X1 U19 ( .A0(data2_i[14]), .A1(select_i), .B0(data1_i[14]), .B1(n4), .Y(
        data_o[14]) );
  AO22X1 U20 ( .A0(data2_i[0]), .A1(select_i), .B0(data1_i[0]), .B1(n2), .Y(
        data_o[0]) );
  AO22X1 U21 ( .A0(data2_i[4]), .A1(select_i), .B0(data1_i[4]), .B1(n6), .Y(
        data_o[4]) );
  AO22X1 U22 ( .A0(data2_i[6]), .A1(select_i), .B0(data1_i[6]), .B1(n6), .Y(
        data_o[6]) );
  AO22X1 U23 ( .A0(data2_i[7]), .A1(select_i), .B0(data1_i[7]), .B1(n6), .Y(
        data_o[7]) );
  AO22X1 U24 ( .A0(data2_i[3]), .A1(select_i), .B0(data1_i[3]), .B1(n6), .Y(
        data_o[3]) );
  AO22X1 U25 ( .A0(data2_i[11]), .A1(select_i), .B0(data1_i[11]), .B1(n3), .Y(
        data_o[11]) );
  AO22X1 U26 ( .A0(data2_i[13]), .A1(select_i), .B0(data1_i[13]), .B1(n4), .Y(
        data_o[13]) );
  AO22X1 U27 ( .A0(data2_i[10]), .A1(select_i), .B0(data1_i[10]), .B1(n2), .Y(
        data_o[10]) );
  AO22X1 U28 ( .A0(data2_i[12]), .A1(select_i), .B0(data1_i[12]), .B1(n3), .Y(
        data_o[12]) );
  AO22X1 U29 ( .A0(data2_i[8]), .A1(select_i), .B0(data1_i[8]), .B1(n6), .Y(
        data_o[8]) );
  AO22X1 U30 ( .A0(data2_i[5]), .A1(select_i), .B0(data1_i[5]), .B1(n6), .Y(
        data_o[5]) );
  AO22X1 U31 ( .A0(data2_i[1]), .A1(select_i), .B0(data1_i[1]), .B1(n5), .Y(
        data_o[1]) );
  AO22X1 U32 ( .A0(data2_i[2]), .A1(select_i), .B0(data1_i[2]), .B1(n5), .Y(
        data_o[2]) );
  AO22X1 U33 ( .A0(data2_i[15]), .A1(select_i), .B0(data1_i[15]), .B1(n5), .Y(
        data_o[15]) );
  AO22X1 U34 ( .A0(data2_i[16]), .A1(select_i), .B0(data1_i[16]), .B1(n5), .Y(
        data_o[16]) );
  AO22X1 U35 ( .A0(data2_i[17]), .A1(select_i), .B0(data1_i[17]), .B1(n5), .Y(
        data_o[17]) );
  AO22X1 U36 ( .A0(data2_i[22]), .A1(select_i), .B0(data1_i[22]), .B1(n5), .Y(
        data_o[22]) );
  AO22X1 U37 ( .A0(data2_i[25]), .A1(select_i), .B0(data1_i[25]), .B1(n5), .Y(
        data_o[25]) );
  AO22X1 U38 ( .A0(data2_i[27]), .A1(select_i), .B0(data1_i[27]), .B1(n5), .Y(
        data_o[27]) );
  AO22X1 U39 ( .A0(select_i), .A1(data2_i[9]), .B0(data1_i[9]), .B1(n6), .Y(
        data_o[9]) );
endmodule


module Mux_WIDTH32_3 ( data1_i, data2_i, select_i, data_o );
  input [31:0] data1_i;
  input [31:0] data2_i;
  output [31:0] data_o;
  input select_i;
  wire   n1, n2, n3, n4, n5, n6, n7;

  CLKBUFX3 U1 ( .A(n7), .Y(n4) );
  CLKBUFX3 U2 ( .A(n4), .Y(n2) );
  CLKBUFX3 U3 ( .A(n7), .Y(n3) );
  CLKBUFX3 U4 ( .A(n7), .Y(n5) );
  CLKBUFX3 U5 ( .A(n7), .Y(n6) );
  AO22X1 U6 ( .A0(data2_i[31]), .A1(n1), .B0(data1_i[31]), .B1(n6), .Y(
        data_o[31]) );
  AO22X1 U7 ( .A0(data2_i[30]), .A1(select_i), .B0(data1_i[30]), .B1(n6), .Y(
        data_o[30]) );
  AO22X1 U8 ( .A0(data2_i[18]), .A1(select_i), .B0(data1_i[18]), .B1(n5), .Y(
        data_o[18]) );
  AO22X1 U9 ( .A0(data2_i[19]), .A1(n1), .B0(data1_i[19]), .B1(n5), .Y(
        data_o[19]) );
  AO22X1 U10 ( .A0(data2_i[20]), .A1(n1), .B0(data1_i[20]), .B1(n5), .Y(
        data_o[20]) );
  AO22X1 U11 ( .A0(data2_i[21]), .A1(select_i), .B0(data1_i[21]), .B1(n5), .Y(
        data_o[21]) );
  AO22X1 U12 ( .A0(data2_i[23]), .A1(n1), .B0(data1_i[23]), .B1(n5), .Y(
        data_o[23]) );
  AO22X1 U13 ( .A0(data2_i[24]), .A1(select_i), .B0(data1_i[24]), .B1(n5), .Y(
        data_o[24]) );
  AO22X1 U14 ( .A0(data2_i[26]), .A1(n1), .B0(data1_i[26]), .B1(n5), .Y(
        data_o[26]) );
  AO22X1 U15 ( .A0(data2_i[28]), .A1(select_i), .B0(data1_i[28]), .B1(n5), .Y(
        data_o[28]) );
  AO22X1 U16 ( .A0(data2_i[29]), .A1(n1), .B0(data1_i[29]), .B1(n5), .Y(
        data_o[29]) );
  CLKINVX1 U17 ( .A(n1), .Y(n7) );
  AO22X1 U18 ( .A0(data2_i[14]), .A1(select_i), .B0(data1_i[14]), .B1(n4), .Y(
        data_o[14]) );
  AO22X1 U19 ( .A0(data2_i[0]), .A1(n1), .B0(data1_i[0]), .B1(n2), .Y(
        data_o[0]) );
  AO22X1 U20 ( .A0(data2_i[4]), .A1(select_i), .B0(data1_i[4]), .B1(n6), .Y(
        data_o[4]) );
  AO22X1 U21 ( .A0(data2_i[6]), .A1(n1), .B0(data1_i[6]), .B1(n6), .Y(
        data_o[6]) );
  AO22X1 U22 ( .A0(data2_i[7]), .A1(select_i), .B0(data1_i[7]), .B1(n6), .Y(
        data_o[7]) );
  AO22X1 U23 ( .A0(data2_i[3]), .A1(n1), .B0(data1_i[3]), .B1(n6), .Y(
        data_o[3]) );
  AO22X1 U24 ( .A0(data2_i[11]), .A1(select_i), .B0(data1_i[11]), .B1(n3), .Y(
        data_o[11]) );
  AO22X1 U25 ( .A0(data2_i[13]), .A1(n1), .B0(data1_i[13]), .B1(n4), .Y(
        data_o[13]) );
  AO22X1 U26 ( .A0(data2_i[10]), .A1(select_i), .B0(data1_i[10]), .B1(n2), .Y(
        data_o[10]) );
  AO22X1 U27 ( .A0(data2_i[12]), .A1(n1), .B0(data1_i[12]), .B1(n3), .Y(
        data_o[12]) );
  AO22X1 U28 ( .A0(data2_i[8]), .A1(select_i), .B0(data1_i[8]), .B1(n6), .Y(
        data_o[8]) );
  AO22X1 U29 ( .A0(data2_i[5]), .A1(n1), .B0(data1_i[5]), .B1(n6), .Y(
        data_o[5]) );
  AO22X1 U30 ( .A0(data2_i[1]), .A1(select_i), .B0(data1_i[1]), .B1(n5), .Y(
        data_o[1]) );
  AO22X1 U31 ( .A0(data2_i[2]), .A1(select_i), .B0(data1_i[2]), .B1(n5), .Y(
        data_o[2]) );
  AO22X1 U32 ( .A0(data2_i[15]), .A1(n1), .B0(data1_i[15]), .B1(n5), .Y(
        data_o[15]) );
  AO22X1 U33 ( .A0(data2_i[16]), .A1(select_i), .B0(data1_i[16]), .B1(n5), .Y(
        data_o[16]) );
  AO22X1 U34 ( .A0(data2_i[17]), .A1(n1), .B0(data1_i[17]), .B1(n5), .Y(
        data_o[17]) );
  AO22X1 U35 ( .A0(data2_i[22]), .A1(n1), .B0(data1_i[22]), .B1(n5), .Y(
        data_o[22]) );
  AO22X1 U36 ( .A0(data2_i[25]), .A1(select_i), .B0(data1_i[25]), .B1(n5), .Y(
        data_o[25]) );
  AO22X1 U37 ( .A0(data2_i[27]), .A1(n1), .B0(data1_i[27]), .B1(n5), .Y(
        data_o[27]) );
  AO22X1 U38 ( .A0(select_i), .A1(data2_i[9]), .B0(data1_i[9]), .B1(n6), .Y(
        data_o[9]) );
  CLKBUFX3 U39 ( .A(select_i), .Y(n1) );
endmodule


module Mux_WIDTH32_2 ( data1_i, data2_i, select_i, data_o );
  input [31:0] data1_i;
  input [31:0] data2_i;
  output [31:0] data_o;
  input select_i;
  wire   n1, n2, n3, n4, n5, n6, n7;

  CLKBUFX3 U1 ( .A(n7), .Y(n4) );
  CLKBUFX3 U2 ( .A(n4), .Y(n2) );
  CLKBUFX3 U3 ( .A(n7), .Y(n3) );
  CLKBUFX3 U4 ( .A(n7), .Y(n5) );
  CLKBUFX3 U5 ( .A(n7), .Y(n6) );
  AO22X1 U6 ( .A0(data2_i[31]), .A1(n1), .B0(data1_i[31]), .B1(n6), .Y(
        data_o[31]) );
  AO22X1 U7 ( .A0(data2_i[30]), .A1(select_i), .B0(data1_i[30]), .B1(n6), .Y(
        data_o[30]) );
  AO22X1 U8 ( .A0(data2_i[18]), .A1(select_i), .B0(data1_i[18]), .B1(n5), .Y(
        data_o[18]) );
  AO22X1 U9 ( .A0(data2_i[19]), .A1(n1), .B0(data1_i[19]), .B1(n5), .Y(
        data_o[19]) );
  AO22X1 U10 ( .A0(data2_i[20]), .A1(n1), .B0(data1_i[20]), .B1(n5), .Y(
        data_o[20]) );
  AO22X1 U11 ( .A0(data2_i[21]), .A1(select_i), .B0(data1_i[21]), .B1(n5), .Y(
        data_o[21]) );
  AO22X1 U12 ( .A0(data2_i[23]), .A1(n1), .B0(data1_i[23]), .B1(n5), .Y(
        data_o[23]) );
  AO22X1 U13 ( .A0(data2_i[24]), .A1(select_i), .B0(data1_i[24]), .B1(n5), .Y(
        data_o[24]) );
  AO22X1 U14 ( .A0(data2_i[26]), .A1(n1), .B0(data1_i[26]), .B1(n5), .Y(
        data_o[26]) );
  AO22X1 U15 ( .A0(data2_i[28]), .A1(select_i), .B0(data1_i[28]), .B1(n5), .Y(
        data_o[28]) );
  AO22X1 U16 ( .A0(data2_i[29]), .A1(n1), .B0(data1_i[29]), .B1(n5), .Y(
        data_o[29]) );
  CLKINVX1 U17 ( .A(n1), .Y(n7) );
  AO22X1 U18 ( .A0(data2_i[14]), .A1(select_i), .B0(data1_i[14]), .B1(n4), .Y(
        data_o[14]) );
  AO22X1 U19 ( .A0(data2_i[0]), .A1(n1), .B0(data1_i[0]), .B1(n2), .Y(
        data_o[0]) );
  AO22X1 U20 ( .A0(data2_i[4]), .A1(select_i), .B0(data1_i[4]), .B1(n6), .Y(
        data_o[4]) );
  AO22X1 U21 ( .A0(data2_i[6]), .A1(n1), .B0(data1_i[6]), .B1(n6), .Y(
        data_o[6]) );
  AO22X1 U22 ( .A0(data2_i[7]), .A1(select_i), .B0(data1_i[7]), .B1(n6), .Y(
        data_o[7]) );
  AO22X1 U23 ( .A0(data2_i[3]), .A1(n1), .B0(data1_i[3]), .B1(n6), .Y(
        data_o[3]) );
  AO22X1 U24 ( .A0(data2_i[11]), .A1(select_i), .B0(data1_i[11]), .B1(n3), .Y(
        data_o[11]) );
  AO22X1 U25 ( .A0(data2_i[13]), .A1(n1), .B0(data1_i[13]), .B1(n4), .Y(
        data_o[13]) );
  AO22X1 U26 ( .A0(data2_i[10]), .A1(select_i), .B0(data1_i[10]), .B1(n2), .Y(
        data_o[10]) );
  AO22X1 U27 ( .A0(data2_i[12]), .A1(n1), .B0(data1_i[12]), .B1(n3), .Y(
        data_o[12]) );
  AO22X1 U28 ( .A0(data2_i[8]), .A1(select_i), .B0(data1_i[8]), .B1(n6), .Y(
        data_o[8]) );
  AO22X1 U29 ( .A0(data2_i[5]), .A1(n1), .B0(data1_i[5]), .B1(n6), .Y(
        data_o[5]) );
  AO22X1 U30 ( .A0(data2_i[1]), .A1(select_i), .B0(data1_i[1]), .B1(n5), .Y(
        data_o[1]) );
  AO22X1 U31 ( .A0(data2_i[2]), .A1(select_i), .B0(data1_i[2]), .B1(n5), .Y(
        data_o[2]) );
  AO22X1 U32 ( .A0(data2_i[15]), .A1(n1), .B0(data1_i[15]), .B1(n5), .Y(
        data_o[15]) );
  AO22X1 U33 ( .A0(data2_i[16]), .A1(select_i), .B0(data1_i[16]), .B1(n5), .Y(
        data_o[16]) );
  AO22X1 U34 ( .A0(data2_i[17]), .A1(n1), .B0(data1_i[17]), .B1(n5), .Y(
        data_o[17]) );
  AO22X1 U35 ( .A0(data2_i[22]), .A1(n1), .B0(data1_i[22]), .B1(n5), .Y(
        data_o[22]) );
  AO22X1 U36 ( .A0(data2_i[25]), .A1(select_i), .B0(data1_i[25]), .B1(n5), .Y(
        data_o[25]) );
  AO22X1 U37 ( .A0(data2_i[27]), .A1(n1), .B0(data1_i[27]), .B1(n5), .Y(
        data_o[27]) );
  AO22X1 U38 ( .A0(select_i), .A1(data2_i[9]), .B0(data1_i[9]), .B1(n6), .Y(
        data_o[9]) );
  CLKBUFX3 U39 ( .A(select_i), .Y(n1) );
endmodule


module Mux_WIDTH5_1 ( data1_i, data2_i, select_i, data_o );
  input [4:0] data1_i;
  input [4:0] data2_i;
  output [4:0] data_o;
  input select_i;
  wire   n1;

  AO22X1 U1 ( .A0(data2_i[2]), .A1(select_i), .B0(data1_i[2]), .B1(n1), .Y(
        data_o[2]) );
  AO22X1 U2 ( .A0(data2_i[0]), .A1(select_i), .B0(data1_i[0]), .B1(n1), .Y(
        data_o[0]) );
  AO22X1 U3 ( .A0(data2_i[1]), .A1(select_i), .B0(data1_i[1]), .B1(n1), .Y(
        data_o[1]) );
  CLKINVX1 U4 ( .A(select_i), .Y(n1) );
  AO22X1 U5 ( .A0(select_i), .A1(data2_i[4]), .B0(data1_i[4]), .B1(n1), .Y(
        data_o[4]) );
  AO22X1 U6 ( .A0(data2_i[3]), .A1(select_i), .B0(data1_i[3]), .B1(n1), .Y(
        data_o[3]) );
endmodule


module Mux_WIDTH32_1 ( data1_i, data2_i, select_i, data_o );
  input [31:0] data1_i;
  input [31:0] data2_i;
  output [31:0] data_o;
  input select_i;
  wire   n1, n2, n3, n4, n5, n6, n7;

  CLKBUFX3 U1 ( .A(n7), .Y(n4) );
  CLKBUFX3 U2 ( .A(n4), .Y(n2) );
  CLKBUFX3 U3 ( .A(n7), .Y(n3) );
  CLKBUFX3 U4 ( .A(n7), .Y(n5) );
  CLKBUFX3 U5 ( .A(n7), .Y(n6) );
  CLKINVX1 U6 ( .A(n1), .Y(n7) );
  CLKBUFX3 U7 ( .A(select_i), .Y(n1) );
  AO22X1 U8 ( .A0(data2_i[1]), .A1(n1), .B0(data1_i[1]), .B1(n5), .Y(data_o[1]) );
  AO22X1 U9 ( .A0(data2_i[2]), .A1(n1), .B0(data1_i[2]), .B1(n5), .Y(data_o[2]) );
  AO22X1 U10 ( .A0(data2_i[15]), .A1(select_i), .B0(data1_i[15]), .B1(n5), .Y(
        data_o[15]) );
  AO22X1 U11 ( .A0(data2_i[16]), .A1(n1), .B0(data1_i[16]), .B1(n5), .Y(
        data_o[16]) );
  AO22X1 U12 ( .A0(data2_i[17]), .A1(select_i), .B0(data1_i[17]), .B1(n5), .Y(
        data_o[17]) );
  AO22X1 U13 ( .A0(data2_i[18]), .A1(n1), .B0(data1_i[18]), .B1(n5), .Y(
        data_o[18]) );
  AO22X1 U14 ( .A0(data2_i[19]), .A1(select_i), .B0(data1_i[19]), .B1(n5), .Y(
        data_o[19]) );
  AO22X1 U15 ( .A0(data2_i[20]), .A1(select_i), .B0(data1_i[20]), .B1(n5), .Y(
        data_o[20]) );
  AO22X1 U16 ( .A0(data2_i[21]), .A1(n1), .B0(data1_i[21]), .B1(n5), .Y(
        data_o[21]) );
  AO22X1 U17 ( .A0(data2_i[22]), .A1(select_i), .B0(data1_i[22]), .B1(n5), .Y(
        data_o[22]) );
  AO22X1 U18 ( .A0(data2_i[23]), .A1(n1), .B0(data1_i[23]), .B1(n5), .Y(
        data_o[23]) );
  AO22X1 U19 ( .A0(data2_i[24]), .A1(select_i), .B0(data1_i[24]), .B1(n5), .Y(
        data_o[24]) );
  AO22X1 U20 ( .A0(data2_i[25]), .A1(n1), .B0(data1_i[25]), .B1(n5), .Y(
        data_o[25]) );
  AO22X1 U21 ( .A0(data2_i[26]), .A1(n1), .B0(data1_i[26]), .B1(n5), .Y(
        data_o[26]) );
  AO22X1 U22 ( .A0(data2_i[27]), .A1(select_i), .B0(data1_i[27]), .B1(n5), .Y(
        data_o[27]) );
  AO22X1 U23 ( .A0(data2_i[28]), .A1(n1), .B0(data1_i[28]), .B1(n5), .Y(
        data_o[28]) );
  AO22X1 U24 ( .A0(data2_i[29]), .A1(select_i), .B0(data1_i[29]), .B1(n5), .Y(
        data_o[29]) );
  AO22X1 U25 ( .A0(data2_i[10]), .A1(n1), .B0(data1_i[10]), .B1(n2), .Y(
        data_o[10]) );
  AO22X1 U26 ( .A0(data2_i[11]), .A1(select_i), .B0(data1_i[11]), .B1(n3), .Y(
        data_o[11]) );
  AO22X1 U27 ( .A0(data2_i[12]), .A1(n1), .B0(data1_i[12]), .B1(n3), .Y(
        data_o[12]) );
  AO22X1 U28 ( .A0(data2_i[13]), .A1(select_i), .B0(data1_i[13]), .B1(n4), .Y(
        data_o[13]) );
  AO22X1 U29 ( .A0(data2_i[14]), .A1(n1), .B0(data1_i[14]), .B1(n4), .Y(
        data_o[14]) );
  AO22X1 U30 ( .A0(data2_i[0]), .A1(select_i), .B0(data1_i[0]), .B1(n2), .Y(
        data_o[0]) );
  AO22X1 U31 ( .A0(data2_i[3]), .A1(n1), .B0(data1_i[3]), .B1(n6), .Y(
        data_o[3]) );
  AO22X1 U32 ( .A0(data2_i[4]), .A1(n1), .B0(data1_i[4]), .B1(n6), .Y(
        data_o[4]) );
  AO22X1 U33 ( .A0(data2_i[5]), .A1(n1), .B0(data1_i[5]), .B1(n6), .Y(
        data_o[5]) );
  AO22X1 U34 ( .A0(data2_i[6]), .A1(n1), .B0(data1_i[6]), .B1(n6), .Y(
        data_o[6]) );
  AO22X1 U35 ( .A0(data2_i[7]), .A1(n1), .B0(data1_i[7]), .B1(n6), .Y(
        data_o[7]) );
  AO22X1 U36 ( .A0(data2_i[8]), .A1(n1), .B0(data1_i[8]), .B1(n6), .Y(
        data_o[8]) );
  AO22X1 U37 ( .A0(n1), .A1(data2_i[9]), .B0(data1_i[9]), .B1(n6), .Y(
        data_o[9]) );
  AO22X1 U38 ( .A0(data2_i[30]), .A1(select_i), .B0(data1_i[30]), .B1(n6), .Y(
        data_o[30]) );
  AO22X1 U39 ( .A0(data2_i[31]), .A1(select_i), .B0(data1_i[31]), .B1(n6), .Y(
        data_o[31]) );
endmodule


module SingleCycle_MIPS ( clk, rst_n, IR_addr, IR, RF_writedata, ReadDataMem, 
        CEN, WEN, A, ReadData2, OEN );
  output [31:0] IR_addr;
  input [31:0] IR;
  output [31:0] RF_writedata;
  input [31:0] ReadDataMem;
  output [6:0] A;
  output [31:0] ReadData2;
  input clk, rst_n;
  output CEN, WEN, OEN;
  wire   RegDST, Jump, Branch, MemRead, MemToReg, MemWrite, ALUSrc, RegWrite,
         JumpRegister, JumpAndLink, ALUresult_1, ALUresult_0, ALUzero, _2_net_,
         n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n15, n16, n17, n18,
         n19, n20, n21;
  wire   [31:0] PCin;
  wire   [1:0] ALUOp;
  wire   [31:0] ALUin1;
  wire   [31:0] ALUin2;
  wire   [31:9] ALUresult;
  wire   [3:0] ALUctrl;
  wire   [31:0] SignExtend;
  wire   [4:0] Reg_W;
  wire   [4:0] MUX_RegDST;
  wire   [31:0] MUX_MemToReg;
  wire   [31:0] PCAdd4;
  wire   [31:0] BranchAddr;
  wire   [31:0] MUX_Branch;
  wire   [31:0] MUX_Jump;

  PC _PC ( .clk(clk), .rst(rst_n), .PCin(PCin), .PCout(IR_addr) );
  mainControl _mainControl ( .opcode_i(IR[31:26]), .funct_i({IR[5:3], n12, n7, 
        IR[0]}), .RegDst_o(RegDST), .Jump_o(Jump), .Branch_o(Branch), 
        .MemRead_o(MemRead), .MemToReg_o(MemToReg), .ALUOp_o(ALUOp), 
        .MemWrite_o(MemWrite), .ALUSrc_o(ALUSrc), .RegWrite_o(RegWrite), 
        .JumpRegister_o(JumpRegister), .JumpAndLink_o(JumpAndLink) );
  ALU _ALU ( .ALUCtrl_i(ALUctrl), .data1_i(ALUin1), .data2_i(ALUin2), .ALU_o({
        ALUresult, A, ALUresult_1, ALUresult_0}), .Zero_o(ALUzero) );
  ALUControl _ALUControl ( .ALUOp_i(ALUOp), .funct_i({IR[5:3], n11, n6, IR[0]}), .ALUctrl_o(ALUctrl) );
  signExtend _signExtend ( .data_i({IR[15:3], n10, n5, IR[0]}), .data_o(
        SignExtend) );
  register_file _regFile ( .clk(clk), .rst(rst_n), .RegWrite_i(RegWrite), 
        .WriteReg_i(Reg_W), .WriteData_i(RF_writedata), .ReadReg1_i({IR[25], 
        n21, IR[23], n20, n19}), .ReadReg2_i({IR[20], n18, n17, n16, n15}), 
        .ReadData1_o(ALUin1), .ReadData2_o(ReadData2) );
  Mux_WIDTH5_0 MUXX_RegDST ( .data1_i({IR[20], n18, n17, n16, n15}), .data2_i(
        IR[15:11]), .select_i(RegDST), .data_o(MUX_RegDST) );
  Mux_WIDTH32_0 MUXX_Src ( .data1_i(ReadData2), .data2_i(SignExtend), 
        .select_i(ALUSrc), .data_o(ALUin2) );
  Mux_WIDTH32_5 MUXX_MemToReg ( .data1_i({ALUresult, A, ALUresult_1, 
        ALUresult_0}), .data2_i(ReadDataMem), .select_i(MemToReg), .data_o(
        MUX_MemToReg) );
  Add_ALU_0 PC_adder ( .data1_i(IR_addr), .data2_i({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b1, 1'b0, 1'b0}), .Add_ALU_o(PCAdd4) );
  Add_ALU_1 branch_adder ( .data1_i(PCAdd4), .data2_i({SignExtend[29:0], 1'b0, 
        1'b0}), .Add_ALU_o(BranchAddr) );
  Mux_WIDTH32_4 MUXX_Branch ( .data1_i(PCAdd4), .data2_i(BranchAddr), 
        .select_i(_2_net_), .data_o(MUX_Branch) );
  Mux_WIDTH32_3 MUXX_Jump ( .data1_i(MUX_Branch), .data2_i({PCAdd4[31:28], 
        IR[25], n21, IR[23], n20, n19, IR[20], n18, n17, n16, n15, IR[15:3], 
        n9, n4, IR[0], 1'b0, 1'b0}), .select_i(Jump), .data_o(MUX_Jump) );
  Mux_WIDTH32_2 MUXX_JumpRegister ( .data1_i(MUX_Jump), .data2_i(ALUin1), 
        .select_i(JumpRegister), .data_o(PCin) );
  Mux_WIDTH5_1 MUXX_JumpAndLink_1 ( .data1_i(MUX_RegDST), .data2_i({1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1}), .select_i(n13), .data_o(Reg_W) );
  Mux_WIDTH32_1 MUXX_JumpAndLink_2 ( .data1_i(MUX_MemToReg), .data2_i(PCAdd4), 
        .select_i(n13), .data_o(RF_writedata) );
  INVXL U7 ( .A(IR[1]), .Y(n3) );
  INVXL U8 ( .A(n3), .Y(n4) );
  INVXL U9 ( .A(n3), .Y(n5) );
  INVXL U10 ( .A(n3), .Y(n6) );
  INVXL U11 ( .A(n3), .Y(n7) );
  INVXL U12 ( .A(IR[2]), .Y(n8) );
  INVXL U13 ( .A(n8), .Y(n9) );
  INVXL U14 ( .A(n8), .Y(n10) );
  INVXL U15 ( .A(n8), .Y(n11) );
  INVXL U16 ( .A(n8), .Y(n12) );
  CLKINVX1 U17 ( .A(MemRead), .Y(OEN) );
  NOR2X1 U18 ( .A(MemWrite), .B(MemToReg), .Y(CEN) );
  CLKINVX1 U19 ( .A(MemWrite), .Y(WEN) );
  AND2X2 U20 ( .A(Branch), .B(ALUzero), .Y(_2_net_) );
  CLKBUFX3 U21 ( .A(JumpAndLink), .Y(n13) );
  CLKBUFX3 U22 ( .A(IR[19]), .Y(n18) );
  CLKBUFX3 U23 ( .A(IR[18]), .Y(n17) );
  CLKBUFX3 U24 ( .A(IR[24]), .Y(n21) );
  CLKBUFX3 U25 ( .A(IR[17]), .Y(n16) );
  CLKBUFX3 U26 ( .A(IR[16]), .Y(n15) );
  CLKBUFX3 U27 ( .A(IR[21]), .Y(n19) );
  CLKBUFX3 U28 ( .A(IR[22]), .Y(n20) );
endmodule

